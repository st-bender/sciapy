netcdf test_v2.2x {
dimensions:
	time = UNLIMITED ; // (2 currently)
	latitude = 18 ;
	altitude = 11 ;
variables:
	double MSIS_Dens(time, latitude, altitude) ;
		MSIS_Dens:_FillValue = NaN ;
		MSIS_Dens:units = "cm^{-3}" ;
		MSIS_Dens:long_name = "MSIS total number density" ;
		MSIS_Dens:model = "NRLMSIS-00" ;
	double MSIS_Temp(time, latitude, altitude) ;
		MSIS_Temp:_FillValue = NaN ;
		MSIS_Temp:units = "K" ;
		MSIS_Temp:long_name = "MSIS temperature" ;
		MSIS_Temp:model = "NRLMSIS-00" ;
	double NO_AKDIAG(time, latitude, altitude) ;
		NO_AKDIAG:_FillValue = NaN ;
		NO_AKDIAG:units = "1" ;
		NO_AKDIAG:long_name = "NO averaging kernel diagonal element" ;
	double NO_APRIORI(time, latitude, altitude) ;
		NO_APRIORI:_FillValue = NaN ;
		NO_APRIORI:units = "cm^{-3}" ;
		NO_APRIORI:long_name = "NO apriori density" ;
	double NO_DENS(time, latitude, altitude) ;
		NO_DENS:_FillValue = NaN ;
		NO_DENS:units = "cm^{-3}" ;
		NO_DENS:long_name = "NO number density" ;
	double NO_ERR(time, latitude, altitude) ;
		NO_ERR:_FillValue = NaN ;
		NO_ERR:units = "cm^{-3}" ;
		NO_ERR:long_name = "NO density measurement error" ;
	double NO_ETOT(time, latitude, altitude) ;
		NO_ETOT:_FillValue = NaN ;
		NO_ETOT:units = "cm^{-3}" ;
		NO_ETOT:long_name = "NO density total error" ;
	double NO_NOEM(time, latitude, altitude) ;
		NO_NOEM:_FillValue = NaN ;
		NO_NOEM:units = "cm^{-3}" ;
		NO_NOEM:long_name = "NOEM NO number density" ;
	double NO_RSTD(time, latitude, altitude) ;
		NO_RSTD:_FillValue = NaN ;
		NO_RSTD:units = "%" ;
		NO_RSTD:long_name = "NO relative standard deviation" ;
	double NO_VMR(time, latitude, altitude) ;
		NO_VMR:_FillValue = NaN ;
		NO_VMR:units = "ppb" ;
		NO_VMR:long_name = "NO volume mixing ratio" ;
	double UTC(time, latitude) ;
		UTC:_FillValue = NaN ;
		UTC:units = "hours" ;
		UTC:long_name = "measurement utc time" ;
	double aacgm_gm_lats(time, latitude) ;
		aacgm_gm_lats:_FillValue = NaN ;
		aacgm_gm_lats:long_name = "geomagnetic_latitude" ;
		aacgm_gm_lats:model = "AACGM" ;
		aacgm_gm_lats:units = "degrees_north" ;
	double aacgm_gm_lons(time, latitude) ;
		aacgm_gm_lons:_FillValue = NaN ;
		aacgm_gm_lons:long_name = "geomagnetic_longitude" ;
		aacgm_gm_lons:model = "AACGM" ;
		aacgm_gm_lons:units = "degrees_east" ;
	double altitude(altitude) ;
		altitude:_FillValue = NaN ;
		altitude:axis = "Z" ;
		altitude:long_name = "altitude" ;
		altitude:standard_name = "altitude" ;
		altitude:units = "km" ;
		altitude:positive = "up" ;
	double app_LST(time, latitude) ;
		app_LST:_FillValue = NaN ;
		app_LST:units = "hours" ;
		app_LST:long_name = "apparent local solar time" ;
	double gm_lats(time, latitude) ;
		gm_lats:_FillValue = NaN ;
		gm_lats:long_name = "geomagnetic_latitude" ;
		gm_lats:model = "IGRF" ;
		gm_lats:units = "degrees_north" ;
	double gm_lons(time, latitude) ;
		gm_lons:_FillValue = NaN ;
		gm_lons:long_name = "geomagnetic_longitude" ;
		gm_lons:model = "IGRF" ;
		gm_lons:units = "degrees_east" ;
	double latitude(latitude) ;
		latitude:_FillValue = NaN ;
		latitude:axis = "Y" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
	double longitude(time, latitude) ;
		longitude:_FillValue = NaN ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
	double mean_LST(time, latitude) ;
		mean_LST:_FillValue = NaN ;
		mean_LST:units = "hours" ;
		mean_LST:long_name = "mean local solar time" ;
	double mean_SZA(time, latitude) ;
		mean_SZA:_FillValue = NaN ;
		mean_SZA:units = "degrees" ;
		mean_SZA:long_name = "solar zenith angle at mean altitude" ;
	int orbit(time) ;
		orbit:axis = "T" ;
		orbit:calendar = "standard" ;
		orbit:long_name = "orbit" ;
		orbit:standard_name = "orbit" ;
		orbit:units = "orbit number" ;
	double time(time) ;
		time:_FillValue = NaN ;
		time:axis = "T" ;
		time:calendar = "standard" ;
		time:long_name = "equatorial crossing time" ;
		time:standard_name = "time" ;
		time:units = "days since 2000-01-01 00:00:00+00:00" ;
	double utc_days(time, latitude) ;
		utc_days:_FillValue = NaN ;
		utc_days:units = "days since 2000-01-01 00:00:00+00:00" ;
		utc_days:long_name = "measurement utc day" ;

// global attributes:
		:version = "2.2" ;
		:L2_data_version = "v6.2" ;
		:software = "sciapy 0.0.7.dev1" ;
		:creation_time = "Thu Mar 12 2020 20:13:13 +00:00 (UTC)" ;
		:author = "The Dude" ;
data:

 MSIS_Dens =
  3.86110274e+15, 1.02654847e+15, 2.28226922e+14, 5.18408033e+13, 
    1.11146245e+13, 1.84965676e+12, 3.72254756e+11, 1.32933828e+11, 
    6.46776553e+10, 3.64086993e+10, 2.23655115e+10,
  4.48113828e+15, 1.11357572e+15, 2.43037321e+14, 5.43718414e+13, 
    1.12215154e+13, 1.84616822e+12, 3.75635363e+11, 1.36184316e+11, 
    6.72284755e+10, 3.83021646e+10, 2.37527564e+10,
  5.01376778e+15, 1.19673156e+15, 2.58974792e+14, 5.49289583e+13, 
    1.05639965e+13, 1.79769467e+12, 3.83402013e+11, 1.38826533e+11, 
    6.86587603e+10, 3.92743264e+10, 2.44453042e+10,
  5.52009214e+15, 1.29797716e+15, 2.84441653e+14, 5.76829125e+13, 
    1.01591547e+13, 1.73531756e+12, 3.95563741e+11, 1.43007135e+11, 
    7.03803408e+10, 4.01864966e+10, 2.49945957e+10,
  5.97435294e+15, 1.42548667e+15, 3.23088046e+14, 6.48680438e+13, 
    1.05693645e+13, 1.70471756e+12, 4.11028867e+11, 1.4863824e+11, 
    7.24772731e+10, 4.11145167e+10, 2.54572759e+10,
  6.33149056e+15, 1.56889284e+15, 3.70966919e+14, 7.63734033e+13, 
    1.1854881e+13, 1.73639401e+12, 4.2854971e+11, 1.55189948e+11, 
    7.48373232e+10, 4.20375371e+10, 2.58303776e+10,
  6.54243245e+15, 1.69750092e+15, 4.13530801e+14, 8.84804226e+13, 
    1.36267103e+13, 1.83668744e+12, 4.47351601e+11, 1.62044253e+11, 
    7.73419356e+10, 4.29771839e+10, 2.61656958e+10,
  6.59972536e+15, 1.77704851e+15, 4.3261869e+14, 9.4720811e+13, 
    1.50801299e+13, 1.97892808e+12, 4.66010571e+11, 1.68289368e+11, 
    7.97073597e+10, 4.38961013e+10, 2.65102522e+10,
  6.56772243e+15, 1.79655135e+15, 4.2259053e+14, 9.14415867e+13, 
    1.53991935e+13, 2.10234217e+12, 4.8100654e+11, 1.72602288e+11, 
    8.13888806e+10, 4.45994693e+10, 2.68159011e+10,
  6.5535397e+15, 1.77991442e+15, 3.96782656e+14, 8.18732138e+13, 
    1.44152264e+13, 2.13738415e+12, 4.87531686e+11, 1.73788654e+11, 
    8.18400659e+10, 4.48254684e+10, 2.69519491e+10,
  6.64898675e+15, 1.77117114e+15, 3.7599658e+14, 7.23357908e+13, 
    1.27118515e+13, 2.0541678e+12, 4.82409633e+11, 1.71544865e+11, 
    8.08837317e+10, 4.442467e+10, 2.67933127e+10,
  6.89030617e+15, 1.80891293e+15, 3.7550426e+14, 6.69040205e+13, 
    1.10421787e+13, 1.88856478e+12, 4.66837637e+11, 1.66844618e+11, 
    7.89138581e+10, 4.3509418e+10, 2.63378457e+10,
  7.24592042e+15, 1.90877133e+15, 4.01469153e+14, 6.65224794e+13, 
    9.84432291e+12, 1.71495133e+12, 4.4664655e+11, 1.61710286e+11, 
    7.68406604e+10, 4.25035026e+10, 2.57897485e+10,
  7.63379066e+15, 2.05813441e+15, 4.51108499e+14, 7.02491653e+13, 
    9.20950954e+12, 1.59671594e+12, 4.29142241e+11, 1.58190812e+11, 
    7.56309069e+10, 4.19280229e+10, 2.54552046e+10,
  7.97234984e+15, 2.22262413e+15, 5.11821872e+14, 7.59565874e+13, 
    9.02223954e+12, 1.55955368e+12, 4.18863103e+11, 1.57067049e+11, 
    7.56260038e+10, 4.19908317e+10, 2.54758167e+10,
  8.23339215e+15, 2.36458244e+15, 5.63845334e+14, 8.0713263e+13, 
    9.04525523e+12, 1.59225131e+12, 4.16001901e+11, 1.5745164e+11, 
    7.6282151e+10, 4.24075664e+10, 2.5704131e+10,
  8.44080576e+15, 2.46205254e+15, 5.91135768e+14, 8.1914021e+13, 
    8.97248013e+12, 1.65689629e+12, 4.17997379e+11, 1.57613428e+11, 
    7.66176454e+10, 4.26675447e+10, 2.58739047e+10,
  8.58672005e+15, 2.51442114e+15, 6.05223396e+14, 8.09442294e+13, 
    8.60822701e+12, 1.67476695e+12, 4.21615096e+11, 1.56421577e+11, 
    7.6118417e+10, 4.26388027e+10, 2.60237827e+10,
  3.92273859e+15, 1.03496634e+15, 2.29285471e+14, 5.19950252e+13, 
    1.11285633e+13, 1.85781222e+12, 3.75196497e+11, 1.34506092e+11, 
    6.5679808e+10, 3.70730206e+10, 2.28159997e+10,
  4.48337551e+15, 1.1194672e+15, 2.43012371e+14, 5.40976756e+13, 
    1.1220681e+13, 1.84901961e+12, 3.77250274e+11, 1.37264311e+11, 
    6.79982168e+10, 3.88421365e+10, 2.41294146e+10,
  4.96737849e+15, 1.19854609e+15, 2.58447354e+14, 5.45820069e+13, 
    1.05615013e+13, 1.79918185e+12, 3.84568078e+11, 1.39685458e+11, 
    6.92876652e+10, 3.97174326e+10, 2.47524402e+10,
  5.49232834e+15, 1.30204905e+15, 2.84553681e+14, 5.75146252e+13, 
    1.01551329e+13, 1.73593208e+12, 3.96258203e+11, 1.43567223e+11, 
    7.07998202e+10, 4.04820469e+10, 2.51974405e+10,
  5.99778854e+15, 1.43382863e+15, 3.24138546e+14, 6.49326056e+13, 
    1.05628647e+13, 1.70398241e+12, 4.10955767e+11, 1.48722827e+11, 
    7.25760168e+10, 4.11910158e+10, 2.55095759e+10,
  6.38727637e+15, 1.57841335e+15, 3.72324426e+14, 7.65665245e+13, 
    1.18457672e+13, 1.73419228e+12, 4.27701684e+11, 1.54805106e+11, 
    7.462656e+10, 4.19056777e+10, 2.5740633e+10,
  6.58849878e+15, 1.70359807e+15, 4.14271615e+14, 8.86195687e+13, 
    1.36182949e+13, 1.83402361e+12, 4.46234642e+11, 1.6147629e+11, 
    7.70047892e+10, 4.27592485e+10, 2.60172667e+10,
  6.6134195e+15, 1.77817507e+15, 4.3246819e+14, 9.47025021e+13, 
    1.50760206e+13, 1.97704506e+12, 4.65224735e+11, 1.67876284e+11, 
    7.94556663e+10, 4.37319872e+10, 2.63985544e+10,
  6.55886741e+15, 1.79490913e+15, 4.2200282e+14, 9.13264444e+13, 
    1.5398744e+13, 2.10159875e+12, 4.807182e+11, 1.72446735e+11, 
    8.12909305e+10, 4.45357106e+10, 2.67734844e+10,
  6.54382846e+15, 1.77826965e+15, 3.96208581e+14, 8.17664425e+13, 
    1.44145634e+13, 2.13685971e+12, 4.87369494e+11, 1.73704382e+11, 
    8.17875025e+10, 4.47932125e+10, 2.69326599e+10,
  6.6499025e+15, 1.7706165e+15, 3.7554906e+14, 7.2270175e+13, 1.27085796e+13, 
    2.05276732e+12, 4.81902059e+11, 1.71290773e+11, 8.07320461e+10, 
    4.4329221e+10, 2.67314873e+10,
  6.89917478e+15, 1.809324e+15, 3.75176566e+14, 6.68664285e+13, 
    1.10381794e+13, 1.88669424e+12, 4.66078336e+11, 1.66466765e+11, 
    7.86895071e+10, 4.33647216e+10, 2.62396361e+10,
  7.25436908e+15, 1.90972812e+15, 4.01299107e+14, 6.65022821e+13, 
    9.84310524e+12, 1.71416114e+12, 4.46285007e+11, 1.61544192e+11, 
    7.67467812e+10, 4.24401082e+10, 2.5742021e+10,
  7.63702555e+15, 2.05897012e+15, 4.51109114e+14, 7.02448592e+13, 
    9.21215106e+12, 1.59770722e+12, 4.29562331e+11, 1.58450309e+11, 
    7.58032875e+10, 4.20381217e+10, 2.55231402e+10,
  7.97279892e+15, 2.22241073e+15, 5.11826185e+14, 7.5957346e+13, 
    9.02583286e+12, 1.56139315e+12, 4.19694608e+11, 1.57566625e+11, 
    7.59591876e+10, 4.22126098e+10, 2.56229098e+10,
  8.23732056e+15, 2.36309557e+15, 5.63623558e+14, 8.06988612e+13, 
    9.04507553e+12, 1.59293403e+12, 4.16388952e+11, 1.57735847e+11, 
    7.64962625e+10, 4.25616089e+10, 2.58126347e+10,
  8.4516058e+15, 2.46078305e+15, 5.90707132e+14, 8.18549177e+13, 
    8.96168581e+12, 1.65374332e+12, 4.1698956e+11, 1.57151071e+11, 
    7.63720795e+10, 4.2530106e+10, 2.57947444e+10,
  8.59247218e+15, 2.51548598e+15, 6.05129212e+14, 8.08859558e+13, 
    8.58799309e+12, 1.6656334e+12, 4.17929413e+11, 1.54389099e+11, 
    7.48245093e+10, 4.17979339e+10, 2.54726294e+10 ;

 MSIS_Temp =
  247.901556, 223.207344, 220.462114, 211.487096, 187.140743, 221.567325, 
    353.185524, 484.777712, 573.763292, 637.953148, 684.302693,
  237.964006, 219.951649, 218.245177, 206.982023, 185.479707, 222.80502, 
    357.303059, 489.551886, 576.361184, 637.141884, 679.7446,
  232.055252, 217.28484, 211.872879, 198.961963, 187.727036, 227.339042, 
    353.743304, 484.396161, 569.669497, 627.492542, 666.74834,
  229.850016, 217.187442, 206.566586, 189.692084, 187.05586, 233.882745, 
    348.779394, 474.649915, 558.765398, 615.064712, 652.79267,
  231.942239, 220.250009, 204.942627, 182.221513, 181.02583, 239.296919, 
    345.015653, 464.605861, 548.215814, 604.78695, 643.109196,
  237.556217, 225.28504, 206.927202, 178.163075, 172.326808, 240.972521, 
    343.197291, 456.636385, 539.907412, 597.845062, 638.201261,
  244.531111, 229.593248, 210.447524, 177.945103, 165.52624, 238.521136, 
    342.551638, 451.401231, 534.050083, 593.473265, 636.240779,
  249.950218, 230.325528, 212.58769, 181.01807, 163.547699, 234.124947, 
    341.875664, 448.720372, 530.751106, 591.362651, 636.189366,
  251.598925, 226.537319, 211.246483, 185.739735, 166.902663, 231.047542, 
    340.888977, 448.456498, 530.678493, 592.428506, 638.844457,
  249.449591, 219.985639, 206.302725, 189.330074, 174.13807, 231.918037, 
    340.715568, 450.914249, 534.707315, 597.958806, 645.745588,
  245.659965, 213.736888, 199.241753, 188.793886, 182.442863, 237.86557, 
    343.183518, 456.667952, 543.310629, 608.622322, 657.89726,
  243.036638, 210.262953, 191.890127, 182.94697, 188.875491, 248.192246, 
    349.631709, 465.987361, 556.146524, 624.082826, 675.318239,
  243.453678, 210.544556, 185.554106, 173.552525, 192.056874, 260.212268, 
    359.909659, 478.162691, 571.667941, 642.594337, 696.439522,
  247.127183, 214.005609, 180.825746, 163.902028, 192.792033, 269.861222, 
    371.999691, 491.208424, 586.944628, 660.581097, 717.264745,
  252.650427, 218.781536, 177.657925, 156.554633, 193.065155, 273.843946, 
    382.62477, 502.4185, 598.578911, 673.702277, 732.435078,
  257.682114, 222.39051, 175.476967, 152.383118, 194.783112, 272.006055, 
    388.644284, 509.595599, 604.636547, 679.535126, 738.603012,
  260.251972, 223.020218, 173.416889, 150.759401, 199.195818, 267.327303, 
    388.259312, 511.901251, 605.593444, 678.83011, 736.120183,
  260.994576, 223.082066, 171.25901, 148.799889, 204.199894, 266.150826, 
    382.467226, 510.922766, 605.572943, 676.965731, 730.862185,
  246.738383, 222.653821, 220.226487, 211.12347, 187.140744, 221.567324, 
    353.172303, 484.130107, 571.670705, 634.122452, 678.721617,
  238.589475, 219.439382, 217.671083, 207.435253, 185.479518, 222.804911, 
    357.326846, 488.816493, 574.028162, 632.943725, 673.723978,
  233.502757, 217.072674, 211.396884, 199.529491, 187.726818, 227.33882, 
    353.773081, 483.722111, 567.570782, 623.780925, 661.508908,
  230.949975, 216.979117, 206.209051, 189.89881, 187.056588, 233.884302, 
    348.791483, 474.154263, 557.237441, 612.381307, 649.027217,
  232.224023, 219.915217, 204.714508, 182.077672, 181.025887, 239.296057, 
    345.009971, 464.366346, 547.468229, 603.463219, 641.238887,
  237.195183, 224.886741, 206.825453, 177.910486, 172.326687, 240.972722, 
    343.184435, 456.603018, 539.80166, 597.654865, 637.928592,
  244.036658, 229.282562, 210.433703, 177.798263, 165.526532, 238.520827, 
    342.543265, 451.45926, 534.238329, 593.818522, 636.744565,
  249.726102, 230.184908, 212.600752, 181.040695, 163.547514, 234.125178, 
    341.876897, 448.78342, 530.958151, 591.748095, 636.759898,
  251.651171, 226.507245, 211.252809, 185.865354, 166.902611, 231.047686, 
    340.895093, 448.503841, 530.83569, 592.723959, 639.285652,
  249.522463, 219.952163, 206.31411, 189.458759, 174.138069, 231.918201, 
    340.721496, 450.967275, 534.884104, 598.292149, 646.244806,
  245.591369, 213.643635, 199.270705, 188.879267, 182.442974, 237.866319, 
    343.1875, 456.740256, 543.551816, 609.07701, 658.57794,
  242.885702, 210.132292, 191.919436, 182.997997, 188.87552, 248.192498, 
    349.634024, 466.035156, 556.305889, 624.383132, 675.767633,
  243.355687, 210.433863, 185.559845, 173.582344, 192.056936, 260.21164, 
    359.910842, 478.093493, 571.436224, 642.155968, 695.78124,
  247.118133, 213.959098, 180.812956, 163.912491, 192.791826, 269.861533, 
    372.001026, 490.97934, 586.173007, 659.112549, 715.045947,
  252.62483, 218.796353, 177.656807, 156.552856, 193.066384, 273.843884, 
    382.622721, 502.114538, 597.545263, 671.715438, 729.405924,
  257.518173, 222.420693, 175.506339, 152.382775, 194.780986, 272.003705, 
    388.64674, 509.37856, 603.893897, 678.103894, 736.413819,
  259.984013, 223.003365, 173.443158, 150.764147, 199.194509, 267.343532, 
    388.260532, 511.996079, 605.908813, 679.426494, 737.021229,
  260.959736, 223.03065, 171.237271, 148.811716, 204.201345, 266.149186, 
    382.470821, 511.935559, 608.961926, 683.383104, 740.511755 ;

 NO_AKDIAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.0643082, 0.382289, 0.544524, 0.615793, 0.598951, 0.61385, 0.594303, 
    0.607201, 0.582212, 0.505521, 0.276377,
  0.140073, 0.604674, 0.755704, 0.793547, 0.783593, 0.76431, 0.74667, 
    0.694106, 0.682025, 0.592799, 0.242383,
  0.0944228, 0.449411, 0.588719, 0.637415, 0.685343, 0.683771, 0.66576, 
    0.611277, 0.59906, 0.555308, 0.160559,
  0.0908882, 0.449847, 0.606411, 0.666852, 0.686014, 0.677353, 0.668386, 
    0.639806, 0.584699, 0.501547, 0.251808,
  0.0622801, 0.405917, 0.565593, 0.628071, 0.634284, 0.656581, 0.641231, 
    0.633894, 0.610713, 0.563, 0.144641,
  0.108064, 0.451313, 0.614014, 0.679094, 0.654779, 0.623497, 0.669455, 
    0.577756, 0.628245, 0.523392, 0.183967,
  0.0738145, 0.354389, 0.547272, 0.659061, 0.649252, 0.624275, 0.639547, 
    0.603924, 0.569379, 0.522482, 0.209727,
  0.0702983, 0.389638, 0.561749, 0.623315, 0.648445, 0.664578, 0.58331, 
    0.586622, 0.583391, 0.535524, 0.138713,
  0.117804, 0.418847, 0.573053, 0.615075, 0.628, 0.618731, 0.68697, 0.607036, 
    0.57524, 0.529491, 0.215394,
  0.0593421, 0.37259, 0.546741, 0.64737, 0.65352, 0.658922, 0.633761, 
    0.608849, 0.571451, 0.533241, 0.179964,
  0.0731159, 0.411016, 0.563692, 0.598699, 0.63155, 0.643268, 0.609911, 
    0.569184, 0.5262, 0.508721, 0.14005,
  0.103461, 0.43735, 0.622881, 0.631503, 0.636967, 0.641602, 0.592245, 
    0.611891, 0.615795, 0.516734, 0.23837,
  0.0704873, 0.378744, 0.57196, 0.624959, 0.579426, 0.589076, 0.630534, 
    0.604201, 0.599238, 0.555138, 0.161288,
  0.104333, 0.48814, 0.657436, 0.665843, 0.669876, 0.655336, 0.634116, 
    0.599581, 0.595017, 0.542386, 0.169438,
  0.0723566, 0.398762, 0.610337, 0.666093, 0.661529, 0.636861, 0.62446, 
    0.596645, 0.560094, 0.519214, 0.244043,
  0.11171, 0.542865, 0.719741, 0.765078, 0.76334, 0.742761, 0.729258, 
    0.688977, 0.666896, 0.568453, 0.226311,
  0.0470979, 0.336084, 0.567294, 0.62423, 0.617833, 0.610806, 0.582861, 
    0.591847, 0.543831, 0.468989, 0.108146,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.0793406, 0.411896, 0.528841, 0.57663, 0.575613, 0.608277, 0.603268, 
    0.625535, 0.577502, 0.519929, 0.211699,
  0.126774, 0.502061, 0.656909, 0.689812, 0.73671, 0.70774, 0.696056, 
    0.641401, 0.64822, 0.559463, 0.185831,
  0.0927776, 0.459485, 0.638727, 0.649431, 0.652188, 0.670033, 0.627428, 
    0.632504, 0.556885, 0.538569, 0.259051,
  0.0705695, 0.405822, 0.579134, 0.623519, 0.689729, 0.663231, 0.647364, 
    0.626248, 0.62435, 0.52277, 0.14215,
  0.13101, 0.474523, 0.607327, 0.656521, 0.641856, 0.631684, 0.668479, 
    0.615606, 0.621096, 0.538259, 0.222135,
  0.0744182, 0.398227, 0.558437, 0.613157, 0.624637, 0.627624, 0.60705, 
    0.613731, 0.621168, 0.541191, 0.18327,
  0.0873967, 0.4157, 0.549083, 0.63421, 0.643806, 0.648493, 0.630492, 
    0.572433, 0.611497, 0.518722, 0.141508,
  0.0935428, 0.401744, 0.560485, 0.612901, 0.663075, 0.621184, 0.619836, 
    0.588949, 0.551109, 0.47594, 0.240829,
  0.066986, 0.380564, 0.559762, 0.573886, 0.638193, 0.591761, 0.596935, 
    0.606763, 0.598474, 0.527489, 0.154741,
  0.0926712, 0.41302, 0.579252, 0.642762, 0.624107, 0.650825, 0.571026, 
    0.551236, 0.544222, 0.481923, 0.149188,
  0.0837544, 0.433505, 0.575692, 0.583052, 0.630573, 0.603605, 0.574065, 
    0.564223, 0.535364, 0.490413, 0.240831,
  0.0695048, 0.356901, 0.550957, 0.589339, 0.589991, 0.605711, 0.624702, 
    0.642811, 0.564361, 0.481757, 0.143507,
  0.105615, 0.424503, 0.616157, 0.629056, 0.661022, 0.608821, 0.629829, 
    0.628363, 0.593661, 0.540915, 0.181519,
  0.0737055, 0.441696, 0.587303, 0.644258, 0.639234, 0.61749, 0.599182, 
    0.575738, 0.574097, 0.470841, 0.229196,
  0.0863047, 0.421714, 0.599808, 0.652477, 0.682645, 0.674216, 0.691614, 
    0.662196, 0.610998, 0.550953, 0.145024,
  0.0945123, 0.462759, 0.656224, 0.688617, 0.634941, 0.637682, 0.645278, 
    0.634688, 0.657122, 0.584334, 0.235111,
  0.044635, 0.328773, 0.546308, 0.52509, 0.439658, 0.426339, 0.286048, 
    0.255994, 0.203114, 0.191932, 0.121528 ;

 NO_APRIORI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NO_DENS =
  70497200, 126345000, 132089000, 145125000, 259042000, 186754000, 83722100, 
    23130600, 42342800, 20060100, 53095600,
  60792500, 154011000, 143110000, 129373000, 340808000, 214653000, 79362300, 
    1502510, 59025500, 5470720, 84244500,
  6027630, 101761000, 53400400, 79550800, 145950000, 215094000, -2173980, 
    -47146900, 82240800, -12974400, 63366200,
  -16141700, 6060170, 19565500, -41321200, 86109400, 48847900, -26519300, 
    -24704500, 11553800, 19233300, 13056700,
  -34216100, -18771800, -981162, -35617100, 22388600, 119954000, -959853, 
    -23126800, 55054800, 35755800, 29990300,
  -44859700, -30435400, 29202600, -15982300, 9007960, 52022900, 679997, 
    -31791200, 29696300, 2521710, 40530600,
  -43489100, -7733180, -21681800, 1500010, -14671900, 42080900, 2385750, 
    -11356700, 11405400, 38906900, 36297500,
  -19673400, -15316200, -74134200, 29664300, 62978400, 48681700, -47769200, 
    -10006300, -38371200, 62239500, 39717000,
  30549200, 57906700, -59022400, 13901500, 80423300, 50716000, 17015600, 
    15381700, 40034300, -25464400, -3122770,
  68772600, 56988100, -20966300, 12352800, 161464000, 28632600, -14112900, 
    47133300, 57565500, -4012270, -2492940,
  85267600, 77004100, 47086500, -23486100, 73809800, -16254900, -5533090, 
    52277200, 44475400, 43635100, 47027900,
  48689300, 28798500, 32484300, 16559100, 51020400, -33988900, 44391000, 
    8979940, 33206000, 56817500, 21112700,
  -1978880, 39887500, 37307300, -5700240, 52851800, 110716000, 43883300, 
    9783560, 126361000, 30787000, -20749500,
  4775850, 31491400, 49221100, -27445900, 48901900, 113439000, -9090030, 
    28883000, 31475400, -52799000, -9711340,
  -39392700, -107628000, -42933200, 7506830, 121787000, 107175000, 22715900, 
    23137600, 65948900, 108271000, 49894800,
  -65644700, -18629300, -16889000, 13105600, 90429100, 56332400, 57074800, 
    94550100, 50035700, -27690400, -29677300,
  -90480400, -27650000, -27173100, 93203500, 110926000, 194236000, -19304500, 
    16312200, 89005200, 16548000, 14264600,
  -51134400, -40383700, -72064800, 41840900, 109347000, 130541000, 67758100, 
    -17655600, 35771300, 6109860, 15970700,
  59287400, 95244800, 154866000, 194345000, 292194000, 177670000, 74172000, 
    22004500, -53775900, -35187200, -4949000,
  54428900, 97670200, 176395000, 196268000, 385126000, 192129000, 66190000, 
    31288800, -87464200, -42200800, 2142880,
  -18419000, -55726400, 57371100, -5088090, 148770000, 51262300, 69835700, 
    52489500, 54808200, 11595000, 23474600,
  -15861400, 24920100, -12844600, 49403000, 127196000, -98028600, 31215800, 
    64875900, 49344000, -42255900, -44441000,
  -29463700, 46025400, 17737300, 17387600, 10447800, -7953760, -10919100, 
    65032700, 37781800, 13893800, -18692000,
  -74232700, -37706300, 18490400, -25450700, 106793000, -21230300, -23635900, 
    38578800, 22446300, 27017800, -13054200,
  -85091400, -79113000, -11541800, 23288000, 46983800, -13367000, 28355200, 
    44263400, 48436800, -30968300, -17436300,
  -70749400, -32335100, -27732200, 52802400, 61154700, 46841600, 43439100, 
    6004750, 23852500, -484931, -12251300,
  -70948600, -212144, -93298800, 37632300, 27313000, -20154900, 29723700, 
    -53764500, 4065700, 88257900, 20565200,
  -58463700, 71164900, 7375580, -49200500, 6211660, -47639600, 69898500, 
    -665151, 45186900, 32076000, 14520300,
  -52342700, 20869400, 36027100, -43658700, 43381900, 71532200, 15338300, 
    60144900, 77476700, 56502700, 3531260,
  -54703400, 6770030, 37268600, -48536900, 75926000, 51021000, -23861100, 
    73885100, 141845000, 46579300, -31061900,
  -57172400, -64608100, 25168200, 57832200, 57799200, 76721400, 57213200, 
    20329600, 99284200, 580596, -9125260,
  -70025000, -10031600, 95165000, 17025300, -37694100, 105713000, 15668100, 
    -17020300, 97954300, 24068300, -6248150,
  -44134400, 48847200, 54807800, 29800800, 50210200, 110862000, 114300000, 
    127088000, 54110500, -34436900, -3168450,
  8561830, 58276600, 70268100, 114509000, 78314200, 36779500, 49633200, 
    37830400, 87060700, 33272300, 31116200,
  -2451020, 112134000, -17223900, -16440700, 201669000, 46032100, 49446100, 
    30002200, 27107700, 41261300, 21038800,
  -7441450, 16082700, -95986200, -13473700, 136707000, 57997100, 97179000, 
    120874000, -716767, -15385500, -8571230 ;

 NO_ERR =
  28233600, 27387400, 22663800, 21380900, 21427900, 20991900, 21525700, 
    21511300, 21753700, 21499200, 19050300,
  33355600, 37205100, 33372400, 32524000, 32739800, 32151600, 33078300, 
    32874600, 33279500, 31523200, 29036600,
  35430800, 32519600, 25695100, 24210700, 24414800, 25026100, 25894600, 
    27396600, 27778000, 23564400, 21547600,
  32701800, 32628600, 28695200, 27917000, 27301600, 27786000, 28356200, 
    29500900, 29615300, 26308600, 18495200,
  31606600, 34221000, 30010100, 28158100, 27749300, 27906000, 28166200, 
    28711500, 29125200, 25006300, 20507600,
  30002700, 33801400, 29570800, 28018900, 27870600, 27693800, 28629900, 
    29343000, 29481600, 26188500, 17494700,
  32372800, 34411200, 30167100, 28059400, 28582500, 29440200, 28150800, 
    30141300, 29521800, 26384800, 19294100,
  30721400, 33975700, 30856200, 28463000, 28527200, 28996400, 28202900, 
    28813700, 29059300, 25600200, 19842500,
  30499300, 33703000, 30026100, 28488600, 28280900, 28119400, 29601200, 
    30117100, 29869600, 26496200, 16949600,
  32842600, 34568000, 30765800, 29480900, 29046900, 29354000, 28226500, 
    29916900, 30168600, 25768000, 19543000,
  29866300, 34016700, 30585600, 28829800, 28324300, 28025700, 28358900, 
    28980800, 29691800, 26320900, 19726700,
  30439200, 33666800, 29323500, 29063000, 28687800, 29047000, 29713100, 
    30124700, 30371500, 27285700, 17609900,
  32095200, 34635800, 29644600, 29010000, 28945600, 29085000, 29706000, 
    29945000, 29638900, 25577600, 20051800,
  30546000, 34028400, 29912700, 27984500, 28245000, 28785600, 28203000, 
    29254200, 29630800, 26443900, 19108800,
  31779000, 33724000, 28650500, 28490400, 28462800, 28777600, 29264600, 
    30064800, 30102100, 26354800, 18944000,
  29791800, 33621100, 29365200, 27789200, 27308700, 27594400, 28080700, 
    28609100, 29096700, 24945600, 20396700,
  29518500, 33496300, 27121600, 25637700, 26022000, 27056900, 27631800, 
    28737300, 28778300, 24501500, 17906800,
  19716900, 30285300, 29265500, 28560600, 28628600, 28695800, 29087700, 
    29413500, 29746900, 27528000, 16565200,
  28916900, 27354600, 22727400, 21450900, 21611000, 21370700, 21453800, 
    21540100, 21837800, 21398300, 18632800,
  34352500, 37171800, 33516400, 32501100, 32896700, 32569200, 32932500, 
    33010800, 33524400, 31235100, 28025700,
  34907000, 33201300, 27739700, 26684700, 25884600, 26973300, 27599600, 
    29259400, 29308900, 26148200, 20734000,
  32413300, 34023100, 29173700, 28321800, 28248400, 27735500, 28420000, 
    27984900, 29198700, 24436000, 20855300,
  30819300, 33245200, 29159300, 28145200, 26868200, 27796600, 28740000, 
    29448700, 29289700, 26673000, 17491100,
  33522900, 34124900, 30151000, 28694500, 28757600, 29359400, 28539600, 
    29689600, 29349200, 25755200, 20070000,
  30920600, 33930200, 30416400, 29046700, 28432800, 28207600, 28058100, 
    28935000, 28783300, 25961800, 19670800,
  31252900, 33423600, 29805800, 28868300, 28555500, 29107300, 29122100, 
    30143300, 29378400, 26692800, 17208400,
  31634200, 34505500, 30702400, 29576400, 28291000, 29202500, 29117600, 
    29668400, 29283200, 25818000, 20733600,
  30281400, 34150300, 29825100, 29226600, 27785000, 27978300, 28529300, 
    29393900, 29772800, 26877100, 18788000,
  31495800, 33712100, 30060900, 28993700, 29368000, 28726500, 30032000, 
    30324700, 30338800, 27222200, 18411400,
  31028600, 34465000, 30195400, 29716600, 29115900, 29111000, 29638100, 
    29612700, 29883800, 25629200, 20449200,
  30276900, 33620200, 29906100, 28622100, 28285600, 28335000, 29139400, 
    29341900, 30138500, 27216500, 18468400,
  32099000, 34254400, 30014200, 29314300, 28649100, 29511900, 29377800, 
    29645300, 30240800, 26754900, 19434900,
  30323600, 34070100, 29854600, 28544500, 28145900, 28434700, 28262600, 
    28767000, 28865500, 25028600, 21108700,
  30143500, 33403800, 28746400, 27551300, 27427300, 28172200, 28382600, 
    28850900, 29867800, 26703700, 17227600,
  28351700, 34067600, 28532400, 26559800, 27467300, 27283700, 27718800, 
    28646700, 28401300, 24328200, 17978400,
  19144700, 31031200, 30265500, 29338200, 28834700, 27961000, 25400400, 
    24835700, 22836900, 22880700, 17756200 ;

 NO_ETOT =
  110302000, 89185000, 84635000, 83783000, 83930900, 83641000, 83962200, 
    83880700, 84177100, 84640700, 86602000,
  90299500, 57740600, 46421600, 42678800, 43547700, 42468400, 44088200, 
    43405100, 45033600, 48764100, 63524800,
  80482000, 41675300, 30519600, 28047300, 28528700, 29612900, 31121400, 
    33966400, 35143600, 39681200, 61501900,
  79883100, 48039400, 39245600, 36389300, 34083600, 34405300, 35640600, 
    38789800, 40042000, 42336600, 64138200,
  80401700, 49223700, 39137700, 35402300, 34506000, 35156900, 35992100, 
    37885500, 41088500, 44584300, 61338200,
  81399300, 51340600, 41363700, 37651200, 37265200, 36255200, 37160100, 
    38109200, 39729100, 41569400, 64788500,
  79884000, 49500900, 39022800, 34838300, 36121800, 38023500, 35417800, 
    40718800, 39089700, 43779400, 63635500,
  81071100, 53622600, 42209700, 36094200, 36867800, 38399100, 37581000, 
    39757000, 41820000, 43825900, 62918200,
  81093700, 52497100, 41891000, 38019900, 36764600, 35951100, 40093100, 
    40396300, 40874000, 42790600, 64949500,
  79724500, 51055100, 41094800, 38311700, 37509100, 38167200, 34873500, 
    39521300, 41781900, 43638400, 62372200,
  81766200, 52987900, 42389300, 37254800, 36874300, 36650900, 37892100, 
    39423600, 42045500, 43535000, 63736200,
  81227500, 51305600, 41232400, 39228900, 37529200, 37110700, 38934200, 
    41034100, 43621300, 44412700, 64942100,
  80156400, 50246400, 38242100, 37515600, 37303400, 37278200, 39858600, 
    39497000, 40048000, 44355600, 61719400,
  80954800, 52384400, 40950800, 38251400, 40333300, 39926000, 37924500, 
    39517400, 40450600, 42447900, 64283000,
  79593500, 47434900, 36540800, 36102800, 35669000, 36353600, 37605800, 
    39771600, 40623900, 43016800, 63962400,
  79991400, 50746800, 38449800, 35269700, 35435200, 36816900, 37960300, 
    39742100, 41968900, 44025200, 61217100,
  76924100, 44958500, 33093100, 30332000, 30756900, 32374400, 33508100, 
    35827300, 37402300, 41636500, 60939500,
  70608100, 51223500, 40021800, 37284700, 37674500, 38141200, 39752400, 
    39592100, 42188500, 45100500, 60791400,
  109709000, 88530700, 84726800, 84034800, 84099100, 83783400, 83858400, 
    83744100, 84278600, 84491000, 87278600,
  89371800, 56283400, 47406000, 44530200, 44845500, 42933200, 43434300, 
    42585300, 45310000, 47629200, 65897100,
  80704800, 46090700, 35553400, 33347800, 31092000, 32791100, 33775200, 
    37326900, 37763300, 41796600, 63155000,
  80262000, 48491100, 37337700, 36344100, 36257300, 35634900, 37903900, 
    37977000, 42088700, 42983000, 60970500,
  80542500, 50980200, 40598200, 37804100, 34392400, 36062700, 36957400, 
    38369300, 38856300, 43678200, 64626800,
  78580400, 48174100, 39264600, 36132800, 36802900, 37833800, 35794800, 
    38879000, 39262300, 43335700, 62115900,
  80489900, 51506800, 41711400, 38752300, 38136800, 38242900, 38985900, 
    39102300, 39171700, 42966800, 63661700,
  80314400, 50973500, 42081600, 37710900, 37045000, 37018500, 37764300, 
    40895300, 39417400, 43839900, 64898000,
  80462300, 51926700, 41570000, 38651500, 35918600, 38381100, 38498500, 
    40480900, 42844100, 46148200, 61732000,
  81437100, 52982400, 41969800, 40900700, 37606500, 39767000, 39678000, 
    39537500, 40846900, 43826100, 64608200,
  80447700, 51017600, 40796900, 37334500, 38108300, 36577200, 40867100, 
    41982400, 43081400, 45833800, 64815500,
  80840100, 50382100, 40702000, 40077400, 37849500, 39163200, 41191300, 
    41947000, 44004600, 45731000, 61820000,
  81216600, 53627600, 42411100, 40114300, 39802800, 39031200, 38440500, 
    37947300, 42293800, 45730000, 64927800,
  79891300, 50642200, 39134400, 37842200, 36048800, 38740800, 37855600, 
    38268800, 41035700, 43511000, 63657800,
  80680100, 49662800, 40119400, 36877900, 37114600, 38546700, 39529800, 
    40660800, 41650300, 46073700, 62130300,
  79697300, 50205000, 39229700, 36133300, 34849700, 35497500, 35050700, 
    36486600, 39783400, 42648200, 64712700,
  77674400, 48882500, 36366500, 33839600, 36492800, 36081800, 36312400, 
    37502400, 37547600, 40843300, 61319000,
  70977000, 52327400, 41489700, 41864800, 45373200, 45660400, 51266200, 
    52686700, 54817500, 55440200, 60973500 ;

 NO_NOEM =
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _ ;

 NO_RSTD =
  40.0492502, 21.6766789, 17.1579768, 14.7327476, 8.27197906, 11.2404018, 
    25.7108935, 92.9993169, 51.3752043, 107.173942, 35.8792442,
  54.8679525, 24.1574303, 23.3194047, 25.1397123, 9.60652332, 14.978407, 
    41.6801176, 2187.97878, 56.3815639, 576.216659, 34.4670572,
  587.806484, 31.95684, 48.1178044, 30.4342634, 16.7281946, 11.6349596, 
    1191.11491, 58.1090167, 33.7764224, 181.622272, 34.0048796,
  202.592044, 538.410639, 146.662237, 67.5609614, 31.7057139, 56.882691, 
    106.926653, 119.415086, 256.325192, 136.786719, 141.652944,
  92.3734733, 182.300046, 3058.62844, 79.0578121, 123.943882, 23.2639178, 
    2934.4285, 124.148174, 52.9021993, 69.936346, 68.3807765,
  66.8811873, 111.05949, 101.260847, 175.312064, 309.399686, 53.2338643, 
    4210.29799, 92.2991268, 99.2770143, 1038.52148, 43.1641772,
  74.4388824, 444.981237, 139.135588, 1870.6142, 194.81117, 69.9609562, 
    1179.95599, 265.405443, 258.840549, 67.8152204, 53.1554515,
  156.157045, 221.828521, 41.6220854, 95.9503511, 45.2968002, 59.5632445, 
    59.0399253, 287.955588, 75.7320595, 41.1317572, 49.959715,
  99.8366569, 58.202246, 50.8723807, 204.931842, 35.1650579, 55.44483, 
    173.965067, 195.798254, 74.6100219, 104.051931, 542.774524,
  47.7553561, 60.6582778, 146.739291, 238.657632, 17.9897067, 102.519506, 
    200.00496, 63.4729586, 52.4074315, 642.22996, 783.933829,
  35.0265517, 44.1751803, 64.9561976, 122.752607, 38.3747145, 172.413857, 
    512.53278, 55.436787, 66.7600516, 60.3204759, 41.9468018,
  62.5172266, 116.9047, 90.2697611, 175.510746, 56.228097, 85.4602532, 
    66.9349643, 335.466607, 91.4638921, 48.0234083, 83.4090382,
  1621.88713, 86.8337198, 79.4605881, 508.92594, 54.7674819, 26.2699158, 
    67.6931771, 306.07468, 23.455734, 83.0792217, 96.6375093,
  639.592952, 108.056168, 60.7721079, 101.962406, 57.758492, 25.3754, 
    310.263002, 101.285185, 94.1395503, 50.0840925, 196.767902,
  80.6723073, 31.3338536, 66.7327383, 379.526378, 23.3709673, 26.851038, 
    128.828706, 129.939147, 45.6445824, 24.3415134, 37.9678844,
  45.3834049, 180.474307, 173.871751, 212.040654, 30.1990178, 48.9849536, 
    49.199822, 30.2581383, 58.1518796, 90.0875394, 68.7282873,
  32.6241926, 121.143942, 99.8104743, 27.5072288, 23.4588825, 13.92991, 
    143.136574, 176.170596, 32.3332794, 148.06321, 125.533138,
  38.558974, 74.9938713, 40.6099788, 68.260004, 26.1814224, 21.9822125, 
    42.9287421, 166.595868, 83.1585657, 450.550422, 103.722442,
  48.7741071, 28.7203081, 14.6755259, 11.0375363, 7.39611354, 12.0283109, 
    28.924392, 97.8895226, 40.6088973, 60.8127387, 376.496262,
  63.1144484, 38.0584866, 19.0007653, 16.5595512, 8.5418019, 16.9517356, 
    49.7544946, 105.503567, 38.3292822, 74.0154215, 1307.85205,
  189.51626, 59.5791223, 48.3513476, 524.454166, 17.3990724, 52.6182009, 
    39.5207609, 55.7433391, 53.4753924, 225.512721, 88.3252537,
  204.353336, 136.528746, 227.128132, 57.3280975, 22.20856, 28.2932736, 
    91.0436382, 43.136049, 59.1737597, 57.8286109, 46.9280619,
  104.600916, 72.2322891, 164.39537, 161.869378, 257.166102, 349.47748, 
    263.208506, 45.2829115, 77.5233049, 191.977717, 93.5753263,
  45.1592088, 90.5018525, 163.062995, 112.745425, 26.9283567, 138.290085, 
    120.74683, 76.9583294, 130.752953, 95.3267846, 153.743623,
  36.3381023, 42.8882737, 263.532551, 124.728186, 60.5161779, 211.024164, 
    98.9522204, 65.3700348, 59.4244459, 83.8334684, 112.815219,
  44.1740849, 103.366311, 107.477229, 54.6723255, 46.6938763, 62.13985, 
    67.041214, 501.990924, 123.166964, 5504.45321, 140.461829,
  44.5874901, 16265.1312, 32.9076044, 78.5931235, 103.580712, 144.890324, 
    97.9608864, 55.1821369, 720.249895, 29.2529054, 100.818859,
  51.7952165, 47.9875613, 404.376334, 59.4030548, 447.303941, 58.7290825, 
    40.8153251, 4419.1319, 65.8881224, 83.7919317, 129.391266,
  60.1722876, 161.538425, 83.4396885, 66.4099023, 67.6964356, 40.1588376, 
    195.797448, 50.4194038, 39.1586116, 48.1785826, 521.383302,
  56.7215201, 509.081939, 81.0210204, 61.2247589, 38.3477333, 57.0568981, 
    124.210954, 40.0793935, 21.0679263, 55.0227247, 65.8337062,
  52.9571961, 52.0371285, 118.824946, 49.4916327, 48.9377016, 36.9323292, 
    50.9312536, 144.330926, 30.3557867, 4687.683, 202.387658,
  45.8393431, 341.464971, 31.5391163, 172.180813, 76.0042022, 27.9170017, 
    187.500718, 174.176131, 30.8723558, 111.1624, 311.050471,
  68.7074028, 69.7483172, 54.4714438, 95.7843414, 56.05614, 25.6487345, 
    24.7266842, 22.6354967, 53.345469, 72.6795966, 666.215342,
  352.068425, 57.3194044, 40.9096019, 24.0603795, 35.0221288, 76.5975611, 
    57.184707, 76.2637984, 34.3068687, 80.2580525, 55.3653724,
  1156.73067, 30.3811511, 165.655862, 161.549082, 13.6199912, 59.2710304, 
    56.0586174, 95.481998, 104.772076, 58.9613027, 85.453543,
  257.271096, 192.947702, 31.5310951, 217.744198, 21.0923362, 48.2110312, 
    26.1377458, 20.5467677, 3186.09813, 148.715999, 207.160466 ;

 NO_VMR =
  18.2583072, 123.077481, 578.761694, 2799.43579, 23306.4104, 100966.841, 
    224905.387, 174000.858, 654674.32, 550969.971, 2373994.44,
  13.5663075, 138.303123, 588.839604, 2379.41178, 30370.9425, 116269.47, 
    211274.837, 11032.9151, 877983.616, 142830.57, 3546725.21,
  1.20221563, 85.0324364, 206.199219, 1448.24884, 13815.794, 119649.907, 
    -5670.23626, -339610.151, 1197819.47, -330353.215, 2592162.46,
  -2.92417221, 4.66893422, 68.785636, -716.350791, 8476.03981, 28149.2569, 
    -67041.7868, -172750.122, 164162.32, 478601.063, 522380.925,
  -5.72716415, -13.1686955, -3.03682545, -549.070049, 2118.25412, 70365.9088, 
    -2335.24474, -155591.186, 759614.672, 869663.634, 1178063.99,
  -7.08517206, -19.3992854, 78.7202268, -209.265259, 759.85242, 29960.3084, 
    1586.74008, -204853.474, 396811.36, 59987.1014, 1569105.98,
  -6.64723715, -4.55562639, -52.4309191, 16.9530158, -1076.70155, 22911.3017, 
    5333.05345, -70083.9418, 147467.217, 905291.982, 1387217.08,
  -2.98094223, -8.61889807, -171.361528, 313.176162, 4176.25051, 24600.035, 
    -102506.687, -59458.8957, -481400.966, 1417882.18, 1498175.11,
  4.6514146, 32.232143, -139.668061, 152.026015, 5222.56573, 24123.5708, 
    35374.9868, 89116.4314, 491889.06, -570957.466, -116452.175,
  10.4939625, 32.0173259, -52.8407673, 150.877185, 11200.934, 13396.0945, 
    -28947.6569, 271210.456, 703390.196, -89508.7133, -92495.7225,
  12.8241495, 43.4763747, 125.231192, -324.681596, 5806.37681, -7913.13153, 
    -11469.6922, 304743.602, 549868.3, 982226.768, 1755210.36,
  7.06634782, 15.9203351, 86.5084726, 247.505305, 4620.50119, -17997.2116, 
    95088.7343, 53822.1736, 420787.943, 1305866.7, 801610.741,
  -0.27310264, 20.8969505, 92.9269403, -85.6889288, 5368.75928, 64559.2666, 
    98250.6191, 60500.5424, 1644454.89, 724340.304, -804563.876,
  0.625619723, 15.3009443, 109.111445, -390.69361, 5309.93532, 71045.1978, 
    -21181.858, 182583.297, 416171.13, -1259277.12, -381507.049,
  -4.9411655, -48.4238422, -83.8830897, 98.8305328, 13498.5332, 68721.5845, 
    54232.2774, 147310.338, 872039.995, 2578443.81, 1958516.21,
  -7.97298353, -7.87847346, -29.9532495, 162.372323, 9997.40722, 35379.0884, 
    137198.411, 600502.48, 655929.327, -652958.95, -1154573.17,
  -10.7194032, -11.2304671, -45.9676126, 1137.82108, 12362.914, 117228.822, 
    -46183.3039, 103494.989, 1161680.18, 387835.768, 551312.225,
  -5.95505614, -16.0608338, -119.071405, 516.910227, 12702.6158, 77945.7702, 
    160710.802, -112871.896, 469942.774, 143293.423, 613696.333,
  15.113778, 92.026954, 675.428755, 3737.76144, 26256.2195, 95633.9926, 
    197688.413, 163594.82, -818758.484, -949132.265, -216909.189,
  12.1401609, 87.2470402, 725.868396, 3628.03018, 34322.8722, 103908.579, 
    175453.815, 227945.631, -1286271.97, -1086469.59, 88807.7907,
  -3.70799206, -46.4949997, 221.9837, -93.2191813, 14086.0656, 28492.006, 
    181595.156, 375769.252, 791023.913, 291937.299, 948375.183,
  -2.88791911, 19.1391407, -45.1394618, 858.96413, 12525.2915, -56470.2969, 
    78776.4133, 451885.178, 696950.923, -1043818.27, -1763710.88,
  -4.91242727, 32.099652, 54.7213536, 267.779182, 989.106675, -4667.74772, 
    -26570.0128, 437274.501, 520582.441, 337301.708, -732744.443,
  -11.6219646, -23.8887362, 49.6620654, -332.399834, 9015.28775, -12242.1834, 
    -55262.5835, 249208.834, 300781.652, 644728.865, -507143.705,
  -12.9151424, -46.4387707, -27.8604654, 262.786203, 3450.05012, -7288.34675, 
    63543.2514, 274117.024, 629010.228, -724247.996, -670181.853,
  -10.6978546, -18.18443, -64.1254099, 557.56077, 4056.4219, 23692.7326, 
    93372.2925, 35768.9, 300198.854, -11088.7026, -464089.807,
  -10.817203, -0.118192056, -221.085727, 412.063562, 1773.71609, -9590.27025, 
    61831.8591, -311774.531, 50014.1894, 1981733.28, 768118.175,
  -8.93417369, 40.0191839, 18.6153969, -601.719954, 430.929458, -22294.2104, 
    143419.933, -3829.21255, 552491.501, 716090.635, 539133.529,
  -7.87119811, 11.7865162, 95.9318071, -604.103975, 3413.59157, 34846.7161, 
    31828.6666, 351127.495, 959677.151, 1274615.23, 132101.142,
  -7.92897727, 3.74174554, 99.3361617, -725.878458, 6878.48942, 27042.5377, 
    -51195.4712, 443842.949, 1802591.04, 1074128.88, -1183777.85,
  -7.88109887, -33.8310461, 62.7168104, 869.6273, 5872.04937, 44757.4025, 
    128198.795, 125845.441, 1293659.47, 13680.361, -354488.872,
  -9.1691457, -4.87214453, 210.95783, 242.370761, -4091.78049, 66165.4392, 
    36474.567, -107417.273, 1292217.04, 572535.095, -244803.342,
  -5.53562186, 21.9793755, 107.082837, 392.335983, 5562.9437, 71001.9765, 
    272340.883, 806566.747, 712362.806, -815796.516, -123656.916,
  1.03939502, 24.6611271, 124.672042, 1418.96674, 8658.21404, 23089.1545, 
    119199.128, 239833.878, 1138103.97, 781744.413, 1205463.93,
  -0.290006427, 45.5684217, -29.158104, -200.851708, 22503.4669, 27835.0936, 
    118578.748, 190913.111, 354942.541, 970166.874, 815623.511,
  -0.866042955, 6.39347631, -158.620999, -166.576507, 15918.3873, 34819.8468, 
    232524.912, 782917.969, -9579.30772, -368092.357, -336487.838 ;

 UTC =
  1.76008492, 1.8267015, 1.88917013, 1.93860666, 1.98716402, 2.03494198, 
    2.08252525, 2.12977343, 2.17699254, 2.22408513, 2.27117682, 2.31814491, 
    2.36510991, 2.41262253, 2.46031892, 2.51196217, 2.56645355, 2.62093096,
  3.43675755, 3.5034732, 3.56589479, 3.61502442, 3.66395003, 3.7115925, 
    3.75923425, 3.80643351, 3.85361659, 3.90071129, 3.94778373, 3.99482065, 
    4.04183767, 4.08921096, 4.13724771, 4.18785429, 4.2489747, 4.31008426 ;

 aacgm_gm_lats =
  86.140811, 70.0870441, 59.4612691, 49.4063312, 39.4062013, 29.3744491, 
    19.3830001, 10.1194714, -6.93261113, -14.9611352, -25.6858764, 
    -36.9770053, -48.097177, -58.7631358, -68.5091646, -75.547919, 
    -76.0241588, -70.1210443,
  83.9774634, 69.5675137, 60.1161466, 50.5023119, 40.4597118, 30.0681583, 
    19.5276305, 9.77635152, -7.33049168, -15.9229081, -26.43431, -37.0302644, 
    -47.0956743, -56.2810885, -64.0424257, -69.3601862, -70.9180774, 
    -69.5146025 ;

 aacgm_gm_lons =
  -151.839646, -141.822335, -149.905851, -155.382611, -159.873691, 
    -163.755572, -167.042116, -169.713557, -171.871721, -173.750411, 
    -175.361754, -136.85086, 176.320347, 168.008116, 153.587717, 123.84859, 
    75.6530435, 25.6785642,
  -145.218143, -159.657872, -171.946591, -215.313339, 175.09346, 171.071156, 
    168.037253, 165.534819, 163.207076, 160.639758, 157.275595, 152.472914, 
    145.5365, 135.427621, 120.201946, 97.0205846, 64.7390013, 19.9088658 ;

 altitude = 60, 70, 80, 90, 100, 110, 120, 130, 140, 150, 160 ;

 app_LST =
  18.2997935, 12.2542101, 11.0561454, 10.5368485, 10.2454059, 10.0551839, 
    9.9170338, 9.80681532, 9.7107011, 9.61886035, 9.52268537, 9.4121868, 
    9.27341846, 9.08286441, 8.79063414, 8.27349072, 7.06746878, 1.00973284,
  18.2997994, 12.2543151, 11.0562033, 10.5365996, 10.2455253, 10.0551544, 
    9.91708281, 9.80678206, 9.71068515, 9.61884652, 9.52263229, 9.41216921, 
    9.2734729, 9.08281285, 8.79089627, 8.27271618, 7.07332325, 1.02221948 ;

 gm_lats =
  78.9724345, 79.7376851, 70.8707707, 60.859081, 50.8127596, 40.8697039, 
    31.051861, 21.3563119, 11.7723644, 2.2860771, -7.11805069, -16.4566919, 
    -25.7483835, -35.0167654, -44.3020714, -53.7095155, -63.7003545, 
    -78.5070738,
  80.5021156, 81.4329049, 70.9878549, 60.5374956, 50.34223, 40.3569915, 
    30.5424094, 20.8674086, 11.3049443, 1.82959494, -7.58389153, -16.9621947, 
    -26.3361574, -35.7471857, -45.2651383, -55.0519109, -65.6896426, 
    -80.4200587 ;

 gm_lons =
  177.243436, 72.3843448, 36.630891, 24.352308, 17.9972526, 13.8774232, 
    10.8029796, 8.27032129, 6.01461259, 3.8728594, 1.7176316, -0.574341705, 
    -3.15289667, -6.23513216, -10.1910279, -15.7571816, -24.670462, 
    -31.8453549,
  167.501097, 31.3844475, 2.89162508, -5.66852831, -10.0613528, -12.9029462, 
    -15.0141476, -16.7422413, -18.2676717, -19.7032883, -21.134657, 
    -22.6435261, -24.3274545, -26.3282199, -28.8866572, -32.4728171, 
    -38.0393905, -27.6953287 ;

 latitude = 85, 75, 65, 55, 45, 35, 25, 15, 5, -5, -15, -25, -35, -45, -55, 
    -65, -75, -85 ;

 longitude =
  251.535, 159.852, 140.944, 132.413, 127.313, 123.743, 120.957, 118.595, 
    116.445, 114.361, 112.212, 109.85, 107.064, 103.493, 98.3941, 89.8623, 
    70.9546, -20.7286,
  226.385, 134.702, 115.794, 107.263, 102.163, 98.5928, 95.8071, 93.4446, 
    91.2954, 89.2114, 87.0621, 84.6996, 81.9139, 78.3434, 73.2441, 64.7123, 
    45.8046, -45.8786 ;

 mean_LST =
  18.5290849, 12.4835015, 11.2854368, 10.76614, 10.4746974, 10.2844753, 
    10.1463252, 10.0361068, 9.93999254, 9.8481518, 9.75197682, 9.64147825, 
    9.50270991, 9.31215586, 9.01992559, 8.50278217, 7.29676022, 1.23902429,
  18.5290909, 12.4836065, 11.2854948, 10.7658911, 10.4748167, 10.2844458, 
    10.1463743, 10.0360735, 9.93997659, 9.84813796, 9.75192373, 9.64146065, 
    9.50276434, 9.3121043, 9.02018771, 8.50200763, 7.3026147, 1.25151092 ;

 mean_SZA =
  106.924155, 91.6278735, 82.3071509, 73.9839657, 66.0787559, 58.5552205, 
    51.5432836, 45.3019004, 40.2307193, 36.8654374, 35.7414797, 37.115569, 
    40.7865058, 46.2647388, 53.0838673, 60.9368626, 69.8730869, 78.2485264,
  106.903579, 91.6073678, 82.2868638, 73.9651901, 66.0595393, 58.5381535, 
    51.5275777, 45.2897645, 40.2224341, 36.862363, 35.7450886, 37.1244434, 
    40.7990836, 46.2815778, 53.1001704, 60.96084, 69.871123, 78.2650263 ;

 orbit = 41454, 41455 ;

 time = 3686.09169, 3686.16155 ;

 utc_days =
  3686.07334, 3686.07611, 3686.07872, 3686.08078, 3686.0828, 3686.08479, 
    3686.08677, 3686.08874, 3686.09071, 3686.09267, 3686.09463, 3686.09659, 
    3686.09855, 3686.10053, 3686.10251, 3686.10467, 3686.10694, 3686.10921,
  3686.1432, 3686.14598, 3686.14858, 3686.15063, 3686.15266, 3686.15465, 
    3686.15663, 3686.1586, 3686.16057, 3686.16253, 3686.16449, 3686.16645, 
    3686.16841, 3686.17038, 3686.17239, 3686.17449, 3686.17704, 3686.17959 ;
}
