netcdf test_v2.2 {
dimensions:
	time = UNLIMITED ; // (2 currently)
	altitude = 11 ;
	latitude = 18 ;
variables:
	int orbit(time) ;
		orbit:axis = "T" ;
		orbit:calendar = "standard" ;
		orbit:long_name = "orbit" ;
		orbit:standard_name = "orbit" ;
		orbit:units = "orbit number" ;
	double time(time) ;
		time:axis = "T" ;
		time:calendar = "standard" ;
		time:long_name = "equatorial crossing time" ;
		time:standard_name = "time" ;
		time:units = "days since 2000-01-01 00:00:00+00:00" ;
	double altitude(altitude) ;
		altitude:axis = "Z" ;
		altitude:long_name = "altitude" ;
		altitude:standard_name = "altitude" ;
		altitude:units = "km" ;
		altitude:positive = "up" ;
	double latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
	double longitude(time, latitude) ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
	double NO_DENS(time, latitude, altitude) ;
		NO_DENS:units = "cm^{-3}" ;
		NO_DENS:long_name = "NO number density" ;
	double NO_ERR(time, latitude, altitude) ;
		NO_ERR:units = "cm^{-3}" ;
		NO_ERR:long_name = "NO density measurement error" ;
	double NO_ETOT(time, latitude, altitude) ;
		NO_ETOT:units = "cm^{-3}" ;
		NO_ETOT:long_name = "NO density total error" ;
	double NO_RSTD(time, latitude, altitude) ;
		NO_RSTD:units = "%" ;
		NO_RSTD:long_name = "NO relative standard deviation" ;
	double NO_AKDIAG(time, latitude, altitude) ;
		NO_AKDIAG:units = "1" ;
		NO_AKDIAG:long_name = "NO averaging kernel diagonal element" ;
	double NO_APRIORI(time, latitude, altitude) ;
		NO_APRIORI:units = "cm^{-3}" ;
		NO_APRIORI:long_name = "NO apriori density" ;
	double MSIS_Temp(time, latitude, altitude) ;
		MSIS_Temp:units = "K" ;
		MSIS_Temp:long_name = "MSIS temperature" ;
		MSIS_Temp:model = "NRLMSIS-00" ;
	double NO_NOEM(time, latitude, altitude) ;
		NO_NOEM:units = "cm^{-3}" ;
		NO_NOEM:long_name = "NOEM NO number density" ;
	double MSIS_Dens(time, latitude, altitude) ;
		MSIS_Dens:units = "cm^{-3}" ;
		MSIS_Dens:long_name = "MSIS total number density" ;
		MSIS_Dens:model = "NRLMSIS-00" ;
	double NO_VMR(time, latitude, altitude) ;
		NO_VMR:units = "ppb" ;
		NO_VMR:long_name = "NO volume mixing ratio" ;
	double app_LST(time, latitude) ;
		app_LST:units = "hours" ;
		app_LST:long_name = "apparent local solar time" ;
	double mean_LST(time, latitude) ;
		mean_LST:units = "hours" ;
		mean_LST:long_name = "mean local solar time" ;
	double mean_SZA(time, latitude) ;
		mean_SZA:units = "degrees" ;
		mean_SZA:long_name = "solar zenith angle at mean altitude" ;
	double UTC(time, latitude) ;
		UTC:units = "hours" ;
		UTC:long_name = "measurement utc time" ;
	double utc_days(time, latitude) ;
		utc_days:long_name = "measurement utc day" ;
		utc_days:units = "days since 2000-01-01 00:00:00+00:00" ;
	double gm_lats(time, latitude) ;
		gm_lats:long_name = "geomagnetic_latitude" ;
		gm_lats:model = "IGRF" ;
		gm_lats:units = "degrees_north" ;
	double gm_lons(time, latitude) ;
		gm_lons:long_name = "geomagnetic_longitude" ;
		gm_lons:model = "IGRF" ;
		gm_lons:units = "degrees_east" ;
	double aacgm_gm_lats(time, latitude) ;
		aacgm_gm_lats:long_name = "geomagnetic_latitude" ;
		aacgm_gm_lats:model = "AACGM" ;
		aacgm_gm_lats:units = "degrees_north" ;
	double aacgm_gm_lons(time, latitude) ;
		aacgm_gm_lons:long_name = "geomagnetic_longitude" ;
		aacgm_gm_lons:model = "AACGM" ;
		aacgm_gm_lons:units = "degrees_east" ;

// global attributes:
		:L2_data_version = "v6.2" ;
		:creation_time = "Sat Feb 22 2020 18:33:02 +00:00 (UTC)" ;
		:author = "The Dude" ;
		:version = "2.2" ;
data:

 orbit = 41454, 41455 ;

 time = 3686.09168913024, 3686.1615490428 ;

 altitude = 60, 70, 80, 90, 100, 110, 120, 130, 140, 150, 160 ;

 latitude = 85, 75, 65, 55, 45, 35, 25, 15, 5, -5, -15, -25, -35, -45, -55, 
    -65, -75, -85 ;

 longitude =
  251.535, 159.852, 140.944, 132.413, 127.313, 123.743, 120.957, 118.595, 
    116.445, 114.361, 112.212, 109.85, 107.064, 103.493, 98.3941, 89.8623, 
    70.9546, -20.7286,
  226.385, 134.702, 115.794, 107.263, 102.163, 98.5928, 95.8071, 93.4446, 
    91.2954, 89.2114, 87.0621, 84.6996, 81.9139, 78.3434, 73.2441, 64.7123, 
    45.8046, -45.8786 ;

 NO_DENS =
  70497200, 126345000, 132089000, 145125000, 259042000, 186754000, 83722100, 
    23130600, 42342800, 20060100, 53095600,
  60792500, 154011000, 143110000, 129373000, 340808000, 214653000, 79362300, 
    1502510, 59025500, 5470720, 84244500,
  6027630, 101761000, 53400400, 79550800, 145950000, 215094000, -2173980, 
    -47146900, 82240800, -12974400, 63366200,
  -16141700, 6060170, 19565500, -41321200, 86109400, 48847900, -26519300, 
    -24704500, 11553800, 19233300, 13056700,
  -34216100, -18771800, -981162, -35617100, 22388600, 119954000, -959853, 
    -23126800, 55054800, 35755800, 29990300,
  -44859700, -30435400, 29202600, -15982300, 9007960, 52022900, 679997, 
    -31791200, 29696300, 2521710, 40530600,
  -43489100, -7733180, -21681800, 1500010, -14671900, 42080900, 2385750, 
    -11356700, 11405400, 38906900, 36297500,
  -19673400, -15316200, -74134200, 29664300, 62978400, 48681700, -47769200, 
    -10006300, -38371200, 62239500, 39717000,
  30549200, 57906700, -59022400, 13901500, 80423300, 50716000, 17015600, 
    15381700, 40034300, -25464400, -3122770,
  68772600, 56988100, -20966300, 12352800, 161464000, 28632600, -14112900, 
    47133300, 57565500, -4012270, -2492940,
  85267600, 77004100, 47086500, -23486100, 73809800, -16254900, -5533090, 
    52277200, 44475400, 43635100, 47027900,
  48689300, 28798500, 32484300, 16559100, 51020400, -33988900, 44391000, 
    8979940, 33206000, 56817500, 21112700,
  -1978880, 39887500, 37307300, -5700240, 52851800, 110716000, 43883300, 
    9783560, 126361000, 30787000, -20749500,
  4775850, 31491400, 49221100, -27445900, 48901900, 113439000, -9090030, 
    28883000, 31475400, -52799000, -9711340,
  -39392700, -107628000, -42933200, 7506830, 121787000, 107175000, 22715900, 
    23137600, 65948900, 108271000, 49894800,
  -65644700, -18629300, -16889000, 13105600, 90429100, 56332400, 57074800, 
    94550100, 50035700, -27690400, -29677300,
  -90480400, -27650000, -27173100, 93203500, 110926000, 194236000, -19304500, 
    16312200, 89005200, 16548000, 14264600,
  -51134400, -40383700, -72064800, 41840900, 109347000, 130541000, 67758100, 
    -17655600, 35771300, 6109860, 15970700,
  59287400, 95244800, 154866000, 194345000, 292194000, 177670000, 74172000, 
    22004500, -53775900, -35187200, -4949000,
  54428900, 97670200, 176395000, 196268000, 385126000, 192129000, 66190000, 
    31288800, -87464200, -42200800, 2142880,
  -18419000, -55726400, 57371100, -5088090, 148770000, 51262300, 69835700, 
    52489500, 54808200, 11595000, 23474600,
  -15861400, 24920100, -12844600, 49403000, 127196000, -98028600, 31215800, 
    64875900, 49344000, -42255900, -44441000,
  -29463700, 46025400, 17737300, 17387600, 10447800, -7953760, -10919100, 
    65032700, 37781800, 13893800, -18692000,
  -74232700, -37706300, 18490400, -25450700, 106793000, -21230300, -23635900, 
    38578800, 22446300, 27017800, -13054200,
  -85091400, -79113000, -11541800, 23288000, 46983800, -13367000, 28355200, 
    44263400, 48436800, -30968300, -17436300,
  -70749400, -32335100, -27732200, 52802400, 61154700, 46841600, 43439100, 
    6004750, 23852500, -484931, -12251300,
  -70948600, -212144, -93298800, 37632300, 27313000, -20154900, 29723700, 
    -53764500, 4065700, 88257900, 20565200,
  -58463700, 71164900, 7375580, -49200500, 6211660, -47639600, 69898500, 
    -665151, 45186900, 32076000, 14520300,
  -52342700, 20869400, 36027100, -43658700, 43381900, 71532200, 15338300, 
    60144900, 77476700, 56502700, 3531260,
  -54703400, 6770030, 37268600, -48536900, 75926000, 51021000, -23861100, 
    73885100, 141845000, 46579300, -31061900,
  -57172400, -64608100, 25168200, 57832200, 57799200, 76721400, 57213200, 
    20329600, 99284200, 580596, -9125260,
  -70025000, -10031600, 95165000, 17025300, -37694100, 105713000, 15668100, 
    -17020300, 97954300, 24068300, -6248150,
  -44134400, 48847200, 54807800, 29800800, 50210200, 110862000, 114300000, 
    127088000, 54110500, -34436900, -3168450,
  8561830, 58276600, 70268100, 114509000, 78314200, 36779500, 49633200, 
    37830400, 87060700, 33272300, 31116200,
  -2451020, 112134000, -17223900, -16440700, 201669000, 46032100, 49446100, 
    30002200, 27107700, 41261300, 21038800,
  -7441450, 16082700, -95986200, -13473700, 136707000, 57997100, 97179000, 
    120874000, -716767, -15385500, -8571230 ;

 NO_ERR =
  28233600, 27387400, 22663800, 21380900, 21427900, 20991900, 21525700, 
    21511300, 21753700, 21499200, 19050300,
  33355600, 37205100, 33372400, 32524000, 32739800, 32151600, 33078300, 
    32874600, 33279500, 31523200, 29036600,
  35430800, 32519600, 25695100, 24210700, 24414800, 25026100, 25894600, 
    27396600, 27778000, 23564400, 21547600,
  32701800, 32628600, 28695200, 27917000, 27301600, 27786000, 28356200, 
    29500900, 29615300, 26308600, 18495200,
  31606600, 34221000, 30010100, 28158100, 27749300, 27906000, 28166200, 
    28711500, 29125200, 25006300, 20507600,
  30002700, 33801400, 29570800, 28018900, 27870600, 27693800, 28629900, 
    29343000, 29481600, 26188500, 17494700,
  32372800, 34411200, 30167100, 28059400, 28582500, 29440200, 28150800, 
    30141300, 29521800, 26384800, 19294100,
  30721400, 33975700, 30856200, 28463000, 28527200, 28996400, 28202900, 
    28813700, 29059300, 25600200, 19842500,
  30499300, 33703000, 30026100, 28488600, 28280900, 28119400, 29601200, 
    30117100, 29869600, 26496200, 16949600,
  32842600, 34568000, 30765800, 29480900, 29046900, 29354000, 28226500, 
    29916900, 30168600, 25768000, 19543000,
  29866300, 34016700, 30585600, 28829800, 28324300, 28025700, 28358900, 
    28980800, 29691800, 26320900, 19726700,
  30439200, 33666800, 29323500, 29063000, 28687800, 29047000, 29713100, 
    30124700, 30371500, 27285700, 17609900,
  32095200, 34635800, 29644600, 29010000, 28945600, 29085000, 29706000, 
    29945000, 29638900, 25577600, 20051800,
  30546000, 34028400, 29912700, 27984500, 28245000, 28785600, 28203000, 
    29254200, 29630800, 26443900, 19108800,
  31779000, 33724000, 28650500, 28490400, 28462800, 28777600, 29264600, 
    30064800, 30102100, 26354800, 18944000,
  29791800, 33621100, 29365200, 27789200, 27308700, 27594400, 28080700, 
    28609100, 29096700, 24945600, 20396700,
  29518500, 33496300, 27121600, 25637700, 26022000, 27056900, 27631800, 
    28737300, 28778300, 24501500, 17906800,
  19716900, 30285300, 29265500, 28560600, 28628600, 28695800, 29087700, 
    29413500, 29746900, 27528000, 16565200,
  28916900, 27354600, 22727400, 21450900, 21611000, 21370700, 21453800, 
    21540100, 21837800, 21398300, 18632800,
  34352500, 37171800, 33516400, 32501100, 32896700, 32569200, 32932500, 
    33010800, 33524400, 31235100, 28025700,
  34907000, 33201300, 27739700, 26684700, 25884600, 26973300, 27599600, 
    29259400, 29308900, 26148200, 20734000,
  32413300, 34023100, 29173700, 28321800, 28248400, 27735500, 28420000, 
    27984900, 29198700, 24436000, 20855300,
  30819300, 33245200, 29159300, 28145200, 26868200, 27796600, 28740000, 
    29448700, 29289700, 26673000, 17491100,
  33522900, 34124900, 30151000, 28694500, 28757600, 29359400, 28539600, 
    29689600, 29349200, 25755200, 20070000,
  30920600, 33930200, 30416400, 29046700, 28432800, 28207600, 28058100, 
    28935000, 28783300, 25961800, 19670800,
  31252900, 33423600, 29805800, 28868300, 28555500, 29107300, 29122100, 
    30143300, 29378400, 26692800, 17208400,
  31634200, 34505500, 30702400, 29576400, 28291000, 29202500, 29117600, 
    29668400, 29283200, 25818000, 20733600,
  30281400, 34150300, 29825100, 29226600, 27785000, 27978300, 28529300, 
    29393900, 29772800, 26877100, 18788000,
  31495800, 33712100, 30060900, 28993700, 29368000, 28726500, 30032000, 
    30324700, 30338800, 27222200, 18411400,
  31028600, 34465000, 30195400, 29716600, 29115900, 29111000, 29638100, 
    29612700, 29883800, 25629200, 20449200,
  30276900, 33620200, 29906100, 28622100, 28285600, 28335000, 29139400, 
    29341900, 30138500, 27216500, 18468400,
  32099000, 34254400, 30014200, 29314300, 28649100, 29511900, 29377800, 
    29645300, 30240800, 26754900, 19434900,
  30323600, 34070100, 29854600, 28544500, 28145900, 28434700, 28262600, 
    28767000, 28865500, 25028600, 21108700,
  30143500, 33403800, 28746400, 27551300, 27427300, 28172200, 28382600, 
    28850900, 29867800, 26703700, 17227600,
  28351700, 34067600, 28532400, 26559800, 27467300, 27283700, 27718800, 
    28646700, 28401300, 24328200, 17978400,
  19144700, 31031200, 30265500, 29338200, 28834700, 27961000, 25400400, 
    24835700, 22836900, 22880700, 17756200 ;

 NO_ETOT =
  110302000, 89185000, 84635000, 83783000, 83930900, 83641000, 83962200, 
    83880700, 84177100, 84640700, 86602000,
  90299500, 57740600, 46421600, 42678800, 43547700, 42468400, 44088200, 
    43405100, 45033600, 48764100, 63524800,
  80482000, 41675300, 30519600, 28047300, 28528700, 29612900, 31121400, 
    33966400, 35143600, 39681200, 61501900,
  79883100, 48039400, 39245600, 36389300, 34083600, 34405300, 35640600, 
    38789800, 40042000, 42336600, 64138200,
  80401700, 49223700, 39137700, 35402300, 34506000, 35156900, 35992100, 
    37885500, 41088500, 44584300, 61338200,
  81399300, 51340600, 41363700, 37651200, 37265200, 36255200, 37160100, 
    38109200, 39729100, 41569400, 64788500,
  79884000, 49500900, 39022800, 34838300, 36121800, 38023500, 35417800, 
    40718800, 39089700, 43779400, 63635500,
  81071100, 53622600, 42209700, 36094200, 36867800, 38399100, 37581000, 
    39757000, 41820000, 43825900, 62918200,
  81093700, 52497100, 41891000, 38019900, 36764600, 35951100, 40093100, 
    40396300, 40874000, 42790600, 64949500,
  79724500, 51055100, 41094800, 38311700, 37509100, 38167200, 34873500, 
    39521300, 41781900, 43638400, 62372200,
  81766200, 52987900, 42389300, 37254800, 36874300, 36650900, 37892100, 
    39423600, 42045500, 43535000, 63736200,
  81227500, 51305600, 41232400, 39228900, 37529200, 37110700, 38934200, 
    41034100, 43621300, 44412700, 64942100,
  80156400, 50246400, 38242100, 37515600, 37303400, 37278200, 39858600, 
    39497000, 40048000, 44355600, 61719400,
  80954800, 52384400, 40950800, 38251400, 40333300, 39926000, 37924500, 
    39517400, 40450600, 42447900, 64283000,
  79593500, 47434900, 36540800, 36102800, 35669000, 36353600, 37605800, 
    39771600, 40623900, 43016800, 63962400,
  79991400, 50746800, 38449800, 35269700, 35435200, 36816900, 37960300, 
    39742100, 41968900, 44025200, 61217100,
  76924100, 44958500, 33093100, 30332000, 30756900, 32374400, 33508100, 
    35827300, 37402300, 41636500, 60939500,
  70608100, 51223500, 40021800, 37284700, 37674500, 38141200, 39752400, 
    39592100, 42188500, 45100500, 60791400,
  109709000, 88530700, 84726800, 84034800, 84099100, 83783400, 83858400, 
    83744100, 84278600, 84491000, 87278600,
  89371800, 56283400, 47406000, 44530200, 44845500, 42933200, 43434300, 
    42585300, 45310000, 47629200, 65897100,
  80704800, 46090700, 35553400, 33347800, 31092000, 32791100, 33775200, 
    37326900, 37763300, 41796600, 63155000,
  80262000, 48491100, 37337700, 36344100, 36257300, 35634900, 37903900, 
    37977000, 42088700, 42983000, 60970500,
  80542500, 50980200, 40598200, 37804100, 34392400, 36062700, 36957400, 
    38369300, 38856300, 43678200, 64626800,
  78580400, 48174100, 39264600, 36132800, 36802900, 37833800, 35794800, 
    38879000, 39262300, 43335700, 62115900,
  80489900, 51506800, 41711400, 38752300, 38136800, 38242900, 38985900, 
    39102300, 39171700, 42966800, 63661700,
  80314400, 50973500, 42081600, 37710900, 37045000, 37018500, 37764300, 
    40895300, 39417400, 43839900, 64898000,
  80462300, 51926700, 41570000, 38651500, 35918600, 38381100, 38498500, 
    40480900, 42844100, 46148200, 61732000,
  81437100, 52982400, 41969800, 40900700, 37606500, 39767000, 39678000, 
    39537500, 40846900, 43826100, 64608200,
  80447700, 51017600, 40796900, 37334500, 38108300, 36577200, 40867100, 
    41982400, 43081400, 45833800, 64815500,
  80840100, 50382100, 40702000, 40077400, 37849500, 39163200, 41191300, 
    41947000, 44004600, 45731000, 61820000,
  81216600, 53627600, 42411100, 40114300, 39802800, 39031200, 38440500, 
    37947300, 42293800, 45730000, 64927800,
  79891300, 50642200, 39134400, 37842200, 36048800, 38740800, 37855600, 
    38268800, 41035700, 43511000, 63657800,
  80680100, 49662800, 40119400, 36877900, 37114600, 38546700, 39529800, 
    40660800, 41650300, 46073700, 62130300,
  79697300, 50205000, 39229700, 36133300, 34849700, 35497500, 35050700, 
    36486600, 39783400, 42648200, 64712700,
  77674400, 48882500, 36366500, 33839600, 36492800, 36081800, 36312400, 
    37502400, 37547600, 40843300, 61319000,
  70977000, 52327400, 41489700, 41864800, 45373200, 45660400, 51266200, 
    52686700, 54817500, 55440200, 60973500 ;

 NO_RSTD =
  40.049250182986, 21.676678934663, 17.1579768186601, 14.7327476313523, 
    8.27197906131052, 11.2404018120094, 25.7108935394597, 92.9993169221724, 
    51.375204285026, 107.173942303378, 35.8792442311604,
  54.8679524612411, 24.1574303134192, 23.3194046537628, 25.1397123047313, 
    9.6065233210488, 14.9784070103842, 41.6801176377197, 2187.97878217117, 
    56.3815639003482, 576.216658867571, 34.4670571966122,
  587.806484472338, 31.9568400467763, 48.117804361016, 30.4342633889288, 
    16.7281945871874, 11.634959599059, 1191.11491366066, 58.1090167115972, 
    33.7764224083423, 181.622271550129, 34.0048795730216,
  202.592044208479, 538.410638645451, 146.66223710102, 67.5609614435205, 
    31.7057138941858, 56.8826909652206, 106.926653418454, 119.415086320306, 
    256.325191711818, 136.786718867797, 141.652944465294,
  92.3734733064259, 182.300045813401, 3058.62844260173, 79.0578121183364, 
    123.943882154311, 23.2639178351701, 2934.42850103089, 124.14817441237, 
    52.9021992632795, 69.9363459914196, 68.3807764510525,
  66.8811873463264, 111.059489936061, 101.260846636943, 175.312063970768, 
    309.399686499496, 53.2338643174448, 4210.29798660876, 92.2991268023856, 
    99.2770143081798, 1038.52147947226, 43.1641771895802,
  74.438882386621, 444.981236696935, 139.135588373659, 1870.61419590536, 
    194.811169650829, 69.9609561582571, 1179.9559886828, 265.405443482702, 
    258.84054921353, 67.8152204364779, 53.1554514773745,
  156.157044537294, 221.828521434821, 41.6220853533187, 95.9503510954245, 
    45.2968001727576, 59.5632445046085, 59.0399253075203, 287.955587979573, 
    75.7320594612626, 41.131757163859, 49.9597149835083,
  99.8366569337331, 58.2022460267983, 50.87238065548, 204.931841887566, 
    35.165057887453, 55.4448300339144, 173.965067349961, 195.798253769089, 
    74.6100219062154, 104.05193132373, 542.774523900255,
  47.7553560574996, 60.6582777807998, 146.739291148176, 238.657632277702, 
    17.9897066838428, 102.519505738214, 200.004960001134, 63.4729586088816, 
    52.4074315345129, 642.22995959893, 783.933829133473,
  35.0265517031088, 44.1751802826083, 64.9561976362652, 122.75260686108, 
    38.3747144688104, 172.413856744735, 512.53278005599, 55.4367869740537, 
    66.7600516240439, 60.320475947116, 41.9468017921277,
  62.5172265775026, 116.904699897564, 90.2697610845855, 175.510746356988, 
    56.2280969964955, 85.4602532003095, 66.9349642945642, 335.466606681114, 
    91.4638920676986, 48.0234082808994, 83.4090381618647,
  1621.88712807244, 86.8337198370417, 79.4605881422671, 508.925939960423, 
    54.7674819022247, 26.2699158206583, 67.6931771311638, 306.074680382192, 
    23.4557339685504, 83.0792217494397, 96.6375093375744,
  639.592952039951, 108.05616771563, 60.7721078968166, 101.962406042433, 
    57.7584920013333, 25.3753999947108, 310.263002432335, 101.285185056954, 
    94.1395502519428, 50.0840925017519, 196.767902266834,
  80.6723073056683, 31.3338536440331, 66.7327383004295, 379.526377978454, 
    23.3709673446263, 26.8510380219268, 128.828705884425, 129.939146670355, 
    45.6445823963705, 24.3415134246474, 37.9678844288383,
  45.3834049054988, 180.474306603039, 173.871750843744, 212.040654376755, 
    30.1990177940508, 48.9849535968643, 49.1998219879877, 30.2581382780135, 
    58.1518795579956, 90.0875393638228, 68.7282872768075,
  32.6241926428265, 121.143942133816, 99.8104743293919, 27.5072288057852, 
    23.4588824982421, 13.929910006384, 143.136574373851, 176.17059624085, 
    32.3332794039, 148.063210055596, 125.533137977931,
  38.5589739979349, 74.993871289654, 40.6099787968606, 68.2600039674099, 
    26.1814224441457, 21.9822124849664, 42.9287420987306, 166.595867600082, 
    83.1585656657712, 450.550421777258, 103.722441721402,
  48.7741071458691, 28.7203080903104, 14.6755259385533, 11.0375363400139, 
    7.39611354100358, 12.0283109134913, 28.924391953837, 97.8895225976505, 
    40.6088972941411, 60.8127387231721, 376.496261871085,
  63.114448390469, 38.0584866213031, 19.0007653278154, 16.5595512258748, 
    8.54180190379252, 16.9517355526755, 49.7544946366521, 105.503566771497, 
    38.3292821520119, 74.015421508597, 1307.85204957814,
  189.5162603833, 59.5791222831548, 48.35134762973, 524.454166494696, 
    17.3990723936277, 52.6182009000767, 39.5207608715886, 55.7433391440193, 
    53.4753923682953, 225.512721000431, 88.3252536784439,
  204.353335771117, 136.528745871806, 227.128131666225, 57.3280974839585, 
    22.2085600176106, 28.2932735956649, 91.0436381575997, 43.1360489796673, 
    59.1737597276265, 57.8286109158721, 46.9280619247992,
  104.600915703052, 72.232289127308, 164.395370208544, 161.869378177552, 
    257.166101954478, 349.477479833437, 263.208506195566, 45.2829115198969, 
    77.5233048716578, 191.977716679382, 93.5753263428204,
  45.1592088122889, 90.501852475581, 163.062994851382, 112.745425469633, 
    26.9283567275009, 138.290085396815, 120.746830033974, 76.9583294451875, 
    130.752952602433, 95.3267845642502, 153.743622742106,
  36.338102322914, 42.8882737350372, 263.532551248505, 124.728186190313, 
    60.5161779166436, 211.024163985936, 98.9522204040176, 65.3700348369081, 
    59.424445875863, 83.8334684177046, 112.815218825095,
  44.1740848685643, 103.366310912909, 107.477228636747, 54.672325500356, 
    46.693876349651, 62.1398500478207, 67.0412140214691, 501.990923851951, 
    123.166963630647, 5504.45321086918, 140.461828540645,
  44.5874900984657, 16265.1312316163, 32.907604385051, 78.5931234604316, 
    103.580712481236, 144.890324437234, 97.9608864306933, 55.1821369119028, 
    720.249895466955, 29.2529054056351, 100.818859043433,
  51.7952165189682, 47.9875612837227, 404.37633379341, 59.4030548470036, 
    447.303941297495, 58.7290825279809, 40.8153250785067, 4419.13189636639, 
    65.8881224425663, 83.791931662302, 129.391266020674,
  60.172287635143, 161.538424679195, 83.4396884567451, 66.4099022646116, 
    67.696435610243, 40.1588375584702, 195.79744821786, 50.419403806474, 
    39.1586115567648, 48.1785826164059, 521.383302277374,
  56.7215200517701, 509.081939075602, 81.0210203764026, 61.224758894779, 
    38.3477333192846, 57.0568981399816, 124.210954230945, 40.0793935448419, 
    21.0679262575346, 55.0227246867171, 65.8337062446277,
  52.957196129601, 52.0371284715074, 118.824945764894, 49.4916326890556, 
    48.9377015598832, 36.9323291806458, 50.9312536267854, 144.330926334015, 
    30.3557867213514, 4687.68300160525, 202.387657995498,
  45.8393430917529, 341.464970692611, 31.5391162717386, 172.180813260266, 
    76.0042022491584, 27.9170016932638, 187.500718019415, 174.176130855508, 
    30.8723557822372, 111.162400335711, 311.050470939398,
  68.7074028422274, 69.7483172013954, 54.471443845584, 95.7843413599635, 
    56.0561399874926, 25.6487344626653, 24.7266841644794, 22.6354966637291, 
    53.345468994003, 72.6795965955124, 666.215341886411,
  352.068424624175, 57.3194043578383, 40.9096019388599, 24.0603795334865, 
    35.0221288093347, 76.5975611413967, 57.18470701063, 76.2637984266621, 
    34.3068686560067, 80.2580524941167, 55.3653723783753,
  1156.73066723242, 30.3811511227638, 165.655861912807, 161.549082459993, 
    13.6199911736558, 59.2710304331108, 56.058617363149, 95.4819979868143, 
    104.772075830852, 58.961302721921, 85.4535429777364,
  257.271096358909, 192.947701567523, 31.5310950949199, 217.744197956018, 
    21.0923361642052, 48.2110312412172, 26.1377458092798, 20.5467677085229, 
    3186.09813230799, 148.715998830067, 207.160465884126 ;

 NO_AKDIAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.0643082, 0.382289, 0.544524, 0.615793, 0.598951, 0.61385, 0.594303, 
    0.607201, 0.582212, 0.505521, 0.276377,
  0.140073, 0.604674, 0.755704, 0.793547, 0.783593, 0.76431, 0.74667, 
    0.694106, 0.682025, 0.592799, 0.242383,
  0.0944228, 0.449411, 0.588719, 0.637415, 0.685343, 0.683771, 0.66576, 
    0.611277, 0.59906, 0.555308, 0.160559,
  0.0908882, 0.449847, 0.606411, 0.666852, 0.686014, 0.677353, 0.668386, 
    0.639806, 0.584699, 0.501547, 0.251808,
  0.0622801, 0.405917, 0.565593, 0.628071, 0.634284, 0.656581, 0.641231, 
    0.633894, 0.610713, 0.563, 0.144641,
  0.108064, 0.451313, 0.614014, 0.679094, 0.654779, 0.623497, 0.669455, 
    0.577756, 0.628245, 0.523392, 0.183967,
  0.0738145, 0.354389, 0.547272, 0.659061, 0.649252, 0.624275, 0.639547, 
    0.603924, 0.569379, 0.522482, 0.209727,
  0.0702983, 0.389638, 0.561749, 0.623315, 0.648445, 0.664578, 0.58331, 
    0.586622, 0.583391, 0.535524, 0.138713,
  0.117804, 0.418847, 0.573053, 0.615075, 0.628, 0.618731, 0.68697, 0.607036, 
    0.57524, 0.529491, 0.215394,
  0.0593421, 0.37259, 0.546741, 0.64737, 0.65352, 0.658922, 0.633761, 
    0.608849, 0.571451, 0.533241, 0.179964,
  0.0731159, 0.411016, 0.563692, 0.598699, 0.63155, 0.643268, 0.609911, 
    0.569184, 0.5262, 0.508721, 0.14005,
  0.103461, 0.43735, 0.622881, 0.631503, 0.636967, 0.641602, 0.592245, 
    0.611891, 0.615795, 0.516734, 0.23837,
  0.0704873, 0.378744, 0.57196, 0.624959, 0.579426, 0.589076, 0.630534, 
    0.604201, 0.599238, 0.555138, 0.161288,
  0.104333, 0.48814, 0.657436, 0.665843, 0.669876, 0.655336, 0.634116, 
    0.599581, 0.595017, 0.542386, 0.169438,
  0.0723566, 0.398762, 0.610337, 0.666093, 0.661529, 0.636861, 0.62446, 
    0.596645, 0.560094, 0.519214, 0.244043,
  0.11171, 0.542865, 0.719741, 0.765078, 0.76334, 0.742761, 0.729258, 
    0.688977, 0.666896, 0.568453, 0.226311,
  0.0470979, 0.336084, 0.567294, 0.62423, 0.617833, 0.610806, 0.582861, 
    0.591847, 0.543831, 0.468989, 0.108146,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.0793406, 0.411896, 0.528841, 0.57663, 0.575613, 0.608277, 0.603268, 
    0.625535, 0.577502, 0.519929, 0.211699,
  0.126774, 0.502061, 0.656909, 0.689812, 0.73671, 0.70774, 0.696056, 
    0.641401, 0.64822, 0.559463, 0.185831,
  0.0927776, 0.459485, 0.638727, 0.649431, 0.652188, 0.670033, 0.627428, 
    0.632504, 0.556885, 0.538569, 0.259051,
  0.0705695, 0.405822, 0.579134, 0.623519, 0.689729, 0.663231, 0.647364, 
    0.626248, 0.62435, 0.52277, 0.14215,
  0.13101, 0.474523, 0.607327, 0.656521, 0.641856, 0.631684, 0.668479, 
    0.615606, 0.621096, 0.538259, 0.222135,
  0.0744182, 0.398227, 0.558437, 0.613157, 0.624637, 0.627624, 0.60705, 
    0.613731, 0.621168, 0.541191, 0.18327,
  0.0873967, 0.4157, 0.549083, 0.63421, 0.643806, 0.648493, 0.630492, 
    0.572433, 0.611497, 0.518722, 0.141508,
  0.0935428, 0.401744, 0.560485, 0.612901, 0.663075, 0.621184, 0.619836, 
    0.588949, 0.551109, 0.47594, 0.240829,
  0.066986, 0.380564, 0.559762, 0.573886, 0.638193, 0.591761, 0.596935, 
    0.606763, 0.598474, 0.527489, 0.154741,
  0.0926712, 0.41302, 0.579252, 0.642762, 0.624107, 0.650825, 0.571026, 
    0.551236, 0.544222, 0.481923, 0.149188,
  0.0837544, 0.433505, 0.575692, 0.583052, 0.630573, 0.603605, 0.574065, 
    0.564223, 0.535364, 0.490413, 0.240831,
  0.0695048, 0.356901, 0.550957, 0.589339, 0.589991, 0.605711, 0.624702, 
    0.642811, 0.564361, 0.481757, 0.143507,
  0.105615, 0.424503, 0.616157, 0.629056, 0.661022, 0.608821, 0.629829, 
    0.628363, 0.593661, 0.540915, 0.181519,
  0.0737055, 0.441696, 0.587303, 0.644258, 0.639234, 0.61749, 0.599182, 
    0.575738, 0.574097, 0.470841, 0.229196,
  0.0863047, 0.421714, 0.599808, 0.652477, 0.682645, 0.674216, 0.691614, 
    0.662196, 0.610998, 0.550953, 0.145024,
  0.0945123, 0.462759, 0.656224, 0.688617, 0.634941, 0.637682, 0.645278, 
    0.634688, 0.657122, 0.584334, 0.235111,
  0.044635, 0.328773, 0.546308, 0.52509, 0.439658, 0.426339, 0.286048, 
    0.255994, 0.203114, 0.191932, 0.121528 ;

 NO_APRIORI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MSIS_Temp =
  247.901556393688, 223.207344458175, 220.462114211774, 211.487096284436, 
    187.140742834012, 221.56732460397, 353.185523533568, 484.777712452079, 
    573.763292159671, 637.953147558771, 684.302692672837,
  237.96400638267, 219.951648695858, 218.245176772046, 206.98202349192, 
    185.47970657412, 222.805019816886, 357.303059108994, 489.551885565957, 
    576.361183863422, 637.141883661985, 679.744600482994,
  232.055252306508, 217.284839602717, 211.872878749806, 198.961962544584, 
    187.727036455933, 227.339042184916, 353.743304277794, 484.396161086029, 
    569.669496829652, 627.492541672734, 666.74833952144,
  229.850016369469, 217.187441624809, 206.566586196982, 189.69208402133, 
    187.055860361653, 233.882745147439, 348.779394243864, 474.649914510322, 
    558.765397787505, 615.064712354544, 652.792670133095,
  231.942238534514, 220.250009054526, 204.942626754507, 182.221512530913, 
    181.025829736024, 239.296919262543, 345.015653197062, 464.605860877205, 
    548.215814309309, 604.786949679837, 643.109196450424,
  237.556217181162, 225.285040151795, 206.927201515215, 178.16307546185, 
    172.326808162925, 240.972520925225, 343.197290627317, 456.636384920481, 
    539.907412371146, 597.845062211664, 638.201261027763,
  244.531110872163, 229.593248127999, 210.44752352874, 177.945102851515, 
    165.526240282558, 238.521135674473, 342.551637644856, 451.401231134709, 
    534.050083019931, 593.473264860079, 636.24077854451,
  249.95021754184, 230.325527610664, 212.587689613133, 181.018070458191, 
    163.547698892451, 234.124946778502, 341.875664183777, 448.720372404209, 
    530.751105856207, 591.362650672138, 636.189365835209,
  251.598924767248, 226.537319408245, 211.246482982128, 185.739734707501, 
    166.902663237777, 231.047542068462, 340.888976749456, 448.456497945425, 
    530.678492988506, 592.42850559097, 638.844457306322,
  249.449590938261, 219.985638819303, 206.302725346411, 189.330073592648, 
    174.138069864152, 231.918036576789, 340.715568409301, 450.91424894411, 
    534.707315264906, 597.958805617404, 645.745587933637,
  245.659965318137, 213.736888054781, 199.241752594822, 188.793886192989, 
    182.442862656617, 237.865570413015, 343.183518026624, 456.667952448564, 
    543.310629057686, 608.622322151889, 657.897259876003,
  243.036637810145, 210.262953460868, 191.890126753427, 182.946969842856, 
    188.875490561054, 248.192245941551, 349.631709464773, 465.987361193653, 
    556.146524228971, 624.082826476831, 675.318238945338,
  243.453678357994, 210.544555924405, 185.554106167986, 173.55252527451, 
    192.056874279348, 260.212268236282, 359.909658547129, 478.162691191277, 
    571.667941052777, 642.594337497561, 696.439521571856,
  247.127183267045, 214.00560940842, 180.825746035795, 163.902028438249, 
    192.792032756718, 269.861222349283, 371.999691443045, 491.208423865143, 
    586.944627826089, 660.581096917501, 717.2647454835,
  252.650426916232, 218.781535966214, 177.657925376966, 156.554633087488, 
    193.065154774096, 273.843946368058, 382.624770132979, 502.418499987263, 
    598.578910700392, 673.70227655245, 732.435077843275,
  257.682114002737, 222.39050957885, 175.476966693651, 152.383117838279, 
    194.78311202014, 272.006055312594, 388.644284461819, 509.595599271293, 
    604.636546962678, 679.535126163175, 738.603012087569,
  260.251972285512, 223.020217913984, 173.416889435931, 150.75940119171, 
    199.195818139701, 267.327302773089, 388.259311582136, 511.901251069673, 
    605.593443506215, 678.830110223093, 736.120182742378,
  260.994576245194, 223.082065729591, 171.259010233374, 148.799888824059, 
    204.19989415483, 266.150826077488, 382.467226125485, 510.922766258183, 
    605.572943467864, 676.965730849155, 730.862185057805,
  246.738383214277, 222.653821153336, 220.226487031598, 211.12346952017, 
    187.140744168711, 221.567323783144, 353.172303066329, 484.130106682471, 
    571.670705292833, 634.122452247152, 678.721616598731,
  238.589475006449, 219.439381815853, 217.671082559476, 207.435253332146, 
    185.479517937317, 222.804911434279, 357.326846244536, 488.816493427453, 
    574.028161523785, 632.943725172536, 673.72397757341,
  233.502757145209, 217.072673963057, 211.396884341483, 199.529490562845, 
    187.726818134487, 227.338819561796, 353.773080810788, 483.722111116357, 
    567.570781989869, 623.780925471117, 661.508908415283,
  230.949975459253, 216.979116602357, 206.209051375463, 189.898809639685, 
    187.056587525831, 233.884302024725, 348.791483141107, 474.154262515255, 
    557.237441118298, 612.381306762807, 649.027217458742,
  232.224023044264, 219.915217411915, 204.714508438306, 182.077671942977, 
    181.025887138166, 239.296057251226, 345.00997074719, 464.366345788335, 
    547.468229003827, 603.463218873175, 641.238887140811,
  237.195183229789, 224.886741035947, 206.825453296091, 177.910485931541, 
    172.326687376642, 240.972721761619, 343.184434519798, 456.603017648865, 
    539.801659825896, 597.654864853644, 637.928591884298,
  244.036658343358, 229.282562380802, 210.433703336318, 177.79826259691, 
    165.526532094275, 238.520827325353, 342.543265220235, 451.459260431864, 
    534.238329252454, 593.818521593795, 636.744565416022,
  249.726102109355, 230.184908397625, 212.600751748499, 181.04069485775, 
    163.547514405192, 234.125178089123, 341.876896879878, 448.783420023169, 
    530.958150954334, 591.748094593739, 636.759897549522,
  251.651171277379, 226.507245061394, 211.25280892207, 185.865353616977, 
    166.902611376366, 231.047686482865, 340.895092577451, 448.503841194781, 
    530.835689890062, 592.723958678621, 639.285651750814,
  249.522462850396, 219.952163495289, 206.314109618351, 189.458759407252, 
    174.138068502821, 231.918200567457, 340.721496413301, 450.967275264711, 
    534.884103819376, 598.292148857427, 646.244805996413,
  245.591368714066, 213.643634594021, 199.270704860035, 188.879267417345, 
    182.442974327195, 237.866318693668, 343.187500009351, 456.740255718488, 
    543.551816397405, 609.077009846534, 658.577939827689,
  242.885702235156, 210.132291657659, 191.919435882384, 182.99799679092, 
    188.875519963315, 248.192498483947, 349.634024292129, 466.035156082091, 
    556.305888561002, 624.383132164104, 675.767632921174,
  243.355686952048, 210.433863363672, 185.559845425901, 173.582343746514, 
    192.056936457041, 260.211640321395, 359.910841772078, 478.093493372493, 
    571.436223876772, 642.155968201683, 695.781240113943,
  247.118133341495, 213.95909843672, 180.812956099283, 163.912490678701, 
    192.791825756422, 269.86153324856, 372.001026063939, 490.979340480486, 
    586.173006703684, 659.112548897507, 715.045947292354,
  252.624829945489, 218.796353029434, 177.656807242618, 156.552856205923, 
    193.066384496572, 273.843884046443, 382.622721467997, 502.114537810082, 
    597.545262737552, 671.715437790629, 729.405924195637,
  257.518173110807, 222.420692840487, 175.50633914542, 152.382774702684, 
    194.780986154965, 272.003705116551, 388.646740341675, 509.378559523929, 
    603.893897045817, 678.10389421548, 736.413818925484,
  259.98401334516, 223.003364950232, 173.443158454026, 150.764147214168, 
    199.194508656405, 267.343532378431, 388.260531805186, 511.996079145251, 
    605.908812941495, 679.426493857144, 737.0212285613,
  260.959735625014, 223.030649607022, 171.23727128861, 148.811715879153, 
    204.201345388273, 266.149185729899, 382.470820636411, 511.935558604883, 
    608.961926220092, 683.383103515632, 740.511755118029 ;

 NO_NOEM =
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN,
  NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN, NaN ;

 MSIS_Dens =
  3.86110274344407e+15, 1.02654847060901e+15, 228226922195677, 
    51840803316275.2, 11114624510587.4, 1849656763081.22, 372254756126.548, 
    132933827548.928, 64677655286.9237, 36408699271.7485, 22365511528.6142,
  4.48113827738136e+15, 1.11357572003217e+15, 243037321177724, 
    54371841372201.3, 11221515416658.7, 1846168219743.07, 375635363336.284, 
    136184316204.194, 67228475461.5814, 38302164578.0856, 23752756420.3594,
  5.01376777646464e+15, 1.19673155643379e+15, 258974792403857, 
    54928958285521.8, 10563996526693.3, 1797694669515.4, 383402013439.744, 
    138826533311.143, 68658760307.2084, 39274326421.6224, 24445304211.5882,
  5.52009213776137e+15, 1.29797716393327e+15, 284441653084743, 
    57682912529455.9, 10159154735624.3, 1735317564764.14, 395563741081.643, 
    143007134894.921, 70380340800.4289, 40186496608.0718, 24994595655.0054,
  5.9743529446319e+15, 1.42548667485988e+15, 323088045529290, 64868043791544, 
    10569364547850.9, 1704717555550.79, 411028867044.136, 148638240094.292, 
    72477273052.9306, 41114516706.5485, 25457275936.5515,
  6.33149056048023e+15, 1.56889284411579e+15, 370966919122182, 
    76373403333680.6, 11854880970540.2, 1736394006981.37, 428549710399.667, 
    155189948481.879, 74837323157.7178, 42037537115.8097, 25830377559.1909,
  6.54243244841113e+15, 1.69750092217633e+15, 413530801244158, 
    88480422635973.6, 13626710262702.3, 1836687437128.42, 447351601014.885, 
    162044252994.999, 77341935589.3249, 42977183918.2745, 26165695795.5833,
  6.59972535871502e+15, 1.77704851317808e+15, 432618690451455, 
    94720810971763, 15080129858229.9, 1978928081399.46, 466010571499.407, 
    168289368361.412, 79707359741.3911, 43896101285.7963, 26510252181.8202,
  6.56772243435538e+15, 1.79655134714063e+15, 422590529721158, 
    91441586735389, 15399193464109.6, 2102342165053.64, 481006539872.125, 
    172602288483.367, 81388880616.6787, 44599469347.0881, 26815901139.2264,
  6.55353969652556e+15, 1.77991441862258e+15, 396782656261552, 
    81873213776042.8, 14415226398829.9, 2137384148958.98, 487531686076.485, 
    173788653626.716, 81840065920.4861, 44825468429.075, 26951949054.6424,
  6.6489867493953e+15, 1.77117113831373e+15, 375996580162403, 
    72335790833941.5, 12711851547373, 2054167802112.6, 482409632526.82, 
    171544864734.066, 80883731664.7118, 44424669969.2959, 26793312735.2721,
  6.89030616902708e+15, 1.80891293202357e+15, 375504260141073, 
    66904020537028.6, 11042178738526.5, 1888564779619.73, 466837636942.606, 
    166844617987.852, 78913858104.0323, 43509418038.135, 26337845691.1934,
  7.24592042440935e+15, 1.9087713299778e+15, 401469152854184, 
    66522479377260.9, 9844322913643.94, 1714951328328.53, 446646549543.086, 
    161710285807.564, 76840660379.7749, 42503502578.5381, 25789748467.7222,
  7.63379066162938e+15, 2.05813441279417e+15, 451108498900586, 
    70249165307827.1, 9209509538475.07, 1596715942368.3, 429142241300.701, 
    158190812060.942, 75630906893.3964, 41928022858.199, 25455204600.2086,
  7.97234984265022e+15, 2.2226241286601e+15, 511821871778146, 75956587399104, 
    9022239536424.65, 1559553680497.73, 418863103375.176, 157067048595.609, 
    75626003809.3794, 41990831748.9926, 25475816705.0782,
  8.23339215364149e+15, 2.36458243982666e+15, 563845334428440, 
    80713262968258.6, 9045255231840.39, 1592251313120.48, 416001901310.577, 
    157451639592.193, 76282151038.0342, 42407566373.2554, 25704131001.9544,
  8.44080576425603e+15, 2.46205253677042e+15, 591135767898401, 
    81914021015258.2, 8972480134261.04, 1656896288429.36, 417997378963.198, 
    157613427854.661, 76617645381.0894, 42667544738.7234, 25873904737.3408,
  8.58672005031909e+15, 2.51442113830815e+15, 605223395797403, 
    80944229448936.9, 8608227005623.84, 1674766951263.96, 421615095561.908, 
    156421577340.042, 76118416956.4174, 42638802712.8544, 26023782658.2236,
  3.9227385867589e+15, 1.03496634307215e+15, 229285470563321, 
    51995025158285.8, 11128563278193, 1857812218446.35, 375196497407.91, 
    134506092394.044, 65679807964.4375, 37073020605.2827, 22815999740.1926,
  4.48337551379152e+15, 1.1194672021933e+15, 243012370916426, 
    54097675636408.1, 11220680986063.2, 1849019605114.52, 377250274196.331, 
    137264311288.052, 67998216811.3568, 38842136499.2498, 24129414570.0956,
  4.96737849094118e+15, 1.1985460868076e+15, 258447354260124, 54582006915500, 
    10561501296863.8, 1799181848074.91, 384568077723.242, 139685457751.978, 
    69287665168.7849, 39717432626.4464, 24752440184.0287,
  5.49232834282129e+15, 1.30204904851335e+15, 284553680973845, 
    57514625235544.7, 10155132911599.8, 1735932080024.51, 396258203427.586, 
    143567222788.164, 70799820190.1314, 40482046933.729, 25197440521.1193,
  5.99778854299742e+15, 1.43382863061779e+15, 324138546273408, 
    64932605577991.8, 10562864717057.2, 1703982406739.95, 410955767330.183, 
    148722827060.1, 72576016781.8096, 41191015832.1595, 25509575938.2106,
  6.3872763686054e+15, 1.57841334656691e+15, 372324425994732, 
    76566524474630.4, 11845767208326.3, 1734192283384.5, 427701683624.967, 
    154805106421.413, 74626560003.375, 41905677664.626, 25740633044.8556,
  6.58849878038732e+15, 1.7035980672785e+15, 414271614503876, 
    88619568723988.5, 13618294919852.1, 1834023608056.99, 446234641636.073, 
    161476289791.541, 77004789223.7461, 42759248477.0326, 26017266689.3982,
  6.61341949658452e+15, 1.77817506826177e+15, 432468190435250, 
    94702502120486.3, 15076020581613.1, 1977045063319.88, 465224734568.917, 
    167876283816.506, 79455666329.9922, 43731987216.0028, 26398554367.644,
  6.5588674059319e+15, 1.79490913304245e+15, 422002819541584, 
    91326444367527.4, 15398743990374, 2101598754145.72, 480718200226.5, 
    172446735436.994, 81290930544.3944, 44535710567.1879, 26773484434.9069,
  6.5438284550531e+15, 1.77826964834706e+15, 396208580554635, 
    81766442487974.1, 14414563423159.2, 2136859709894.06, 487369494313.892, 
    173704382337.392, 81787502532.5487, 44793212549.8525, 26932659917.6758,
  6.64990250388346e+15, 1.77061649808801e+15, 375549060067325, 
    72270175037043.5, 12708579554581.3, 2052767316632.52, 481902059205.831, 
    171290773076.701, 80732046065.7674, 44329220976.7017, 26731487312.9853,
  6.89917478108848e+15, 1.80932399836562e+15, 375176565806834, 
    66866428505487.3, 11038179369289.5, 1886694235271.49, 466078335732.942, 
    166466765342.173, 78689507058.1563, 43364721561.1047, 26239636090.2357,
  7.25436908197895e+15, 1.90972812034084e+15, 401299106617741, 
    66502282098610.4, 9843105244696.29, 1714161139316.96, 446285006593.455, 
    161544191523.226, 76746781182.3047, 42440108243.2257, 25742021032.5335,
  7.63702555084608e+15, 2.05897012040537e+15, 451109114329898, 
    70244859155306, 9212151058973.97, 1597707222020.2, 429562330647.202, 
    158450308789.823, 75803287495.1679, 42038121707.4724, 25523140155.6313,
  7.97279891618536e+15, 2.22241072819558e+15, 511826185429660, 
    75957346040082.5, 9025832857927.76, 1561393154451.63, 419694608024.821, 
    157566624808.808, 75959187569.0563, 42212609790.0176, 25622909785.788,
  8.23732055736368e+15, 2.36309556575199e+15, 563623558356425, 
    80698861151253.5, 9045075534602.74, 1592934030216.45, 416388951720.593, 
    157735847251.447, 76496262534.1177, 42561608936.3709, 25812634724.8602,
  8.45160580184895e+15, 2.4607830549149e+15, 590707132436446, 
    81854917678193.8, 8961685805856.06, 1653743318927.76, 416989559606.986, 
    157151071429.54, 76372079527.5914, 42530106026.3227, 25794744410.1946,
  8.59247217941316e+15, 2.51548597687405e+15, 605129211695736, 
    80885955786637.5, 8587993087301.61, 1665633403153.85, 417929413061.809, 
    154389099234.833, 74824509348.9898, 41797933892.241, 25472629447.2677 ;

 NO_VMR =
  18.2583071946739, 123.077481110117, 578.761693533902, 2799.43578641341, 
    23306.4103742997, 100966.840836404, 224905.387028926, 174000.857618325, 
    654674.320090276, 550969.971497052, 2373994.43925394,
  13.5663075399506, 138.303123199876, 588.839604166593, 2379.41178255082, 
    30370.942546143, 116269.469761468, 211274.836573232, 11032.9151100421, 
    877983.616239087, 142830.570028151, 3546725.20987042,
  1.20221563278111, 85.0324364331491, 206.199219253451, 1448.24883782601, 
    13815.7940161388, 119649.90698781, -5670.23626322626, -339610.151427845, 
    1197819.4717181, -330353.214991282, 2592162.4640679,
  -2.92417220531144, 4.66893422195181, 68.7856359566681, -716.350790693851, 
    8476.03981245086, 28149.2569382476, -67041.786811614, -172750.122000224, 
    164162.319599475, 478601.063127678, 522380.925069506,
  -5.72716414934006, -13.1686955276837, -3.03682545230864, -549.070049259647, 
    2118.25412006934, 70365.9087743969, -2335.24474060098, -155591.185588103, 
    759614.672033717, 869663.633776947, 1178063.98747244,
  -7.08517205727264, -19.3992853713046, 78.7202267768296, -209.265258615912, 
    759.852420482759, 29960.3084270251, 1586.74007588485, -204853.47350774, 
    396811.360254238, 59987.1013625968, 1569105.98411205,
  -6.64723714656948, -4.55562639110997, -52.4309191353283, 16.9530157667911, 
    -1076.70154550497, 22911.3016996467, 5333.05345188788, -70083.9418251412, 
    147467.217016149, 905291.981763753, 1387217.07550108,
  -2.98094222572778, -8.61889806970347, -171.361528376497, 313.176161560137, 
    4176.25050925074, 24600.0349671997, -102506.687447671, -59458.8956951269, 
    -481400.966290874, 1417882.18490691, 1498175.11080625,
  4.65141459696879, 32.2321430401439, -139.668061276587, 152.02601459911, 
    5222.56572640899, 24123.5707693214, 35374.9868027232, 89116.4313935631, 
    491889.060233566, -570957.465924705, -116452.17454326,
  10.4939625278322, 32.0173258914894, -52.8407672793525, 150.877184738222, 
    11200.9340354936, 13396.0944802298, -28947.6569483649, 271210.456013075, 
    703390.195896583, -89508.7132518962, -92495.7224780223,
  12.8241494852963, 43.4763746620853, 125.231192208349, -324.681595780381, 
    5806.37680710277, -7913.131528633, -11469.6922012485, 304743.602095241, 
    549868.299652202, 982226.767923282, 1755210.35657864,
  7.0663478233907, 15.9203350753781, 86.5084726010724, 247.505304869312, 
    4620.50118985922, -17997.2116216441, 95088.7342561404, 53822.1736385516, 
    420787.942673193, 1305866.69649777, 801610.740967301,
  -0.273102640395241, 20.8969505008565, 92.9269403010652, -85.6889288156702, 
    5368.759280209, 64559.2665932441, 98250.6190742816, 60500.5423813452, 
    1644454.89374346, 724340.30449871, -804563.87645539,
  0.625619723108916, 15.3009442941321, 109.111444630191, -390.69361009108, 
    5309.93532236433, 71045.197827576, -21181.8579603088, 182583.296866022, 
    416171.130201643, -1259277.12304887, -381507.049443256,
  -4.94116550044734, -48.423842165739, -83.8830897375363, 98.8305327694138, 
    13498.5332087804, 68721.5844765247, 54232.2773645053, 147310.337889973, 
    872039.995214196, 2578443.80523845, 1958516.21078959,
  -7.9729835255043, -7.87847346162549, -29.9532495327288, 162.372322937234, 
    9997.40722425152, 35379.088423925, 137198.411401945, 600502.479649556, 
    655929.327098449, -652958.949737402, -1154573.1694934,
  -10.7194031620955, -11.2304670948532, -45.9676126460855, 1137.82108172469, 
    12362.9139702894, 117228.821958509, -46183.3039429169, 103494.989113757, 
    1161680.17898874, 387835.76841209, 551312.22537948,
  -5.95505614487802, -16.0608337977832, -119.071404873653, 516.910226767864, 
    12702.6157568292, 77945.7702467079, 160710.801660684, -112871.895938109, 
    469942.773776829, 143293.423156041, 613696.333455706,
  15.1137779611731, 92.0269539560862, 675.428755339433, 3737.76143791383, 
    26256.2194863528, 95633.992626328, 197688.412638248, 163594.820192505, 
    -818758.484024757, -949132.264528401, -216909.189005725,
  12.1401608748963, 87.2470402068423, 725.868396472145, 3628.03018227848, 
    34322.8722461989, 103908.57915652, 175453.815483652, 227945.630633295, 
    -1286271.96567002, -1086469.58698616, 88807.7907474699,
  -3.70799205931057, -46.4949997445911, 221.983700178477, -93.2191813297929, 
    14086.0655903321, 28492.0059941965, 181595.155826371, 375769.252180846, 
    791023.912647181, 291937.298894775, 948375.183435321,
  -2.88791911370913, 19.1391407477723, -45.1394617565346, 858.964129517937, 
    12525.2915060038, -56470.2969246445, 78776.4132830238, 451885.177828685, 
    696950.922579856, -1043818.26514788, -1763710.88018847,
  -4.91242727028109, 32.0996519508535, 54.7213535814365, 267.779181895226, 
    989.106675117083, -4667.74772353259, -26570.0128043878, 437274.501067142, 
    520582.441353679, 337301.708134921, -732744.442529184,
  -11.6219646240559, -23.8887361678816, 49.6620654167385, -332.399833669254, 
    9015.28774978253, -12242.1834091929, -55262.5834896766, 249208.833557338, 
    300781.651988044, 644728.865053211, -507143.704556596,
  -12.915142407448, -46.4387706933614, -27.8604654432388, 262.786203265466, 
    3450.05011835287, -7288.34674825222, 63543.251362195, 274117.023973874, 
    629010.227653003, -724247.995533273, -670181.853003996,
  -10.6978545722887, -18.1844299681969, -64.1254099453868, 557.560769965946, 
    4056.42189654376, 23692.7325881703, 93372.292512029, 35768.8999511293, 
    300198.854301174, -11088.7025921052, -464089.806940948,
  -10.8172029725488, -0.118192055572421, -221.085726634123, 412.063562318876, 
    1773.71609120028, -9590.27024556491, 61831.859051717, -311774.53063264, 
    50014.1894399849, 1981733.28495234, 768118.174905443,
  -8.93417368770643, 40.0191838544561, 18.6153969449002, -601.719953845812, 
    430.929457774629, -22294.2104151338, 143419.932547074, -3829.21254518528, 
    552491.500544562, 716090.634586682, 539133.529491099,
  -7.87119810695458, 11.7865161781423, 95.9318071347094, -604.103974808722, 
    3413.59156730946, 34846.716147715, 31828.6666491472, 351127.494608645, 
    959677.151460828, 1274615.22569269, 132101.141947483,
  -7.92897726695503, 3.74174553928175, 99.33616168124, -725.87845776774, 
    6878.48941930059, 27042.5377075784, -51195.4711700485, 443842.948759946, 
    1802591.03536089, 1074128.88456728, -1183777.85016457,
  -7.88109887350861, -33.8310460593045, 62.7168104412803, 869.62729962027, 
    5872.04937498191, 44757.4024636744, 128198.794839009, 125845.440856208, 
    1293659.4665014, 13680.3609612064, -354488.87204572,
  -9.16914570126614, -4.87214452535376, 210.95783032751, 242.370761429792, 
    -4091.78049281774, 66165.4391637114, 36474.5669770289, -107417.272519024, 
    1292217.04277989, 572535.094871325, -244803.341669597,
  -5.53562186428708, 21.979375540389, 107.082837025993, 392.335982674726, 
    5562.94369620398, 71001.9764618063, 272340.882666856, 806566.746950437, 
    712362.806024049, -815796.516048235, -123656.915880702,
  1.03939502419221, 24.6611270591823, 124.672042107161, 1418.96674087353, 
    8658.21404148612, 23089.154542704, 119199.128110645, 239833.878342788, 
    1138103.96895104, 781744.413133952, 1205463.9261614,
  -0.290006426880888, 45.5684217168335, -29.1581039980978, -200.851707708452, 
    22503.4669111272, 27835.0935560217, 118578.748222385, 190913.111358912, 
    354942.541406204, 970166.873660334, 815623.510953846,
  -0.866042955347483, 6.39347630949057, -158.620998862409, -166.576507243621, 
    15918.3872891255, 34819.8468463609, 232524.912013378, 782917.968943814, 
    -9579.30771930517, -368092.356901307, -336487.837572629 ;

 app_LST =
  18.2997934720493, 12.2542100510242, 11.0561453513778, 10.5368485464038, 
    10.2454059085678, 10.0551838679824, 9.9170338019505, 9.80681531502381, 
    9.71070109906263, 9.61886035442492, 9.52268537241684, 9.41218680139767, 
    9.27341846234462, 9.08286441414821, 8.790634143296, 8.27349072360098, 
    7.06746877645805, 1.00973284387693,
  18.299799435297, 12.2543150862601, 11.0562033467433, 10.536599642101, 
    10.2455252556644, 10.055154386791, 9.91708280640596, 9.80678206104737, 
    9.71068515011109, 9.61884651594307, 9.52263228525139, 9.41216920554647, 
    9.27347289545712, 9.08281285089891, 8.79089626870463, 8.2727161805631, 
    7.07332325493774, 1.02221947748644 ;

 mean_LST =
  18.5290849168666, 12.4835014958415, 11.2854367961951, 10.7661399912211, 
    10.4746973533851, 10.2844753127997, 10.1463252467678, 10.0361067598411, 
    9.93999254387992, 9.84815179924221, 9.75197681723413, 9.64147824621496, 
    9.50270990716191, 9.3121558589655, 9.01992558811329, 8.50278216841827, 
    7.29676022127534, 1.23902428869422,
  18.5290908801143, 12.4836065310774, 11.2854947915606, 10.7658910869183, 
    10.4748167004817, 10.2844458316083, 10.1463742512233, 10.0360735058647, 
    9.93997659492839, 9.84813796076036, 9.75192373006868, 9.64146065036376, 
    9.50276434027441, 9.3121042957162, 9.02018771352192, 8.50200762538039, 
    7.30261469975503, 1.25151092230373 ;

 mean_SZA =
  106.924154742655, 91.6278735385579, 82.3071509394994, 73.9839657007906, 
    66.0787558513993, 58.5552205442921, 51.5432836401244, 45.3019003910965, 
    40.2307193236288, 36.8654374456471, 35.7414797489146, 37.1155689610858, 
    40.7865057961226, 46.2647388498017, 53.0838672864313, 60.9368625822346, 
    69.8730869289302, 78.2485264372941,
  106.903579043886, 91.6073677620432, 82.286863786175, 73.9651901149983, 
    66.0595393439007, 58.5381535114787, 51.5275776865588, 45.2897645471775, 
    40.2224341184907, 36.8623629594848, 35.7450886132391, 37.1244433831562, 
    40.7990836166126, 46.2815777517464, 53.1001703523131, 60.9608400147367, 
    69.8711230332547, 78.2650263028253 ;

 UTC =
  1.7600849168666, 1.82670149584149, 1.88917012952841, 1.93860665788775, 
    1.98716402005175, 2.03494197946638, 2.08252524676779, 2.12977342650777, 
    2.17699254387992, 2.22408513257554, 2.27117681723413, 2.31814491288162, 
    2.36510990716191, 2.41262252563217, 2.46031892144662, 2.51196216841827, 
    2.56645355460868, 2.62093095536089,
  3.43675754678096, 3.50347319774405, 3.56589479156058, 3.61502442025161, 
    3.66395003381507, 3.71159249827499, 3.75923425122325, 3.80643350586466, 
    3.85361659492839, 3.90071129409369, 3.94778373006868, 3.99482065036376, 
    4.04183767360775, 4.08921096238287, 4.13724771352192, 4.18785429204706, 
    4.24897469975503, 4.31008425563707 ;

 utc_days =
  3686.07333660683, 3686.0761125755, 3686.07871544724, 3686.08077525147, 
    3686.08279855087, 3686.08478920406, 3686.08677193404, 3686.08874052955, 
    3686.09070805424, 3686.09267020624, 3686.09463235825, 3686.09658938824, 
    3686.09854620537, 3686.10052597527, 3686.10251323778, 3686.104665134, 
    3686.10693551561, 3686.10920589723,
  3686.1431979665, 3686.14597806292, 3686.14857899132, 3686.15062599445, 
    3686.1526646118, 3686.1546496816, 3686.15663475139, 3686.15860141238, 
    3686.16056731832, 3686.16252967437, 3686.16449093751, 3686.16645090986, 
    3686.1684098577, 3686.17038383887, 3686.17238528982, 3686.17449397081, 
    3686.17704056711, 3686.17958716341 ;

 gm_lats =
  78.9724344966206, 79.7376850848464, 70.8707706591498, 60.8590810306038, 
    50.8127595658507, 40.8697038681856, 31.0518610288899, 21.3563118781732, 
    11.7723643577302, 2.28607710440003, -7.11805068719162, -16.4566918757602, 
    -25.7483834914115, -35.0167653513888, -44.3020714408483, 
    -53.7095155021783, -63.7003545138594, -78.5070738199646,
  80.5021155597976, 81.4329049438286, 70.9878548849182, 60.5374955597333, 
    50.3422299545729, 40.3569915268545, 30.5424094388205, 20.8674085962378, 
    11.3049443072648, 1.82959494360535, -7.5838915257135, -16.9621946642614, 
    -26.3361573890536, -35.7471856642415, -45.2651382809906, 
    -55.0519108536856, -65.6896426232229, -80.4200587144977 ;

 gm_lons =
  177.243436423979, 72.3843447831355, 36.6308910367747, 24.3523080471894, 
    17.9972525809882, 13.8774232179713, 10.802979619409, 8.27032128928681, 
    6.01461259125558, 3.87285940202976, 1.71763160378014, -0.574341704888147, 
    -3.15289667042224, -6.2351321568916, -10.1910278715936, 
    -15.7571815580906, -24.6704619803908, -31.8453549074452,
  167.501097150302, 31.3844474889351, 2.89162508487009, -5.66852830600422, 
    -10.0613528357414, -12.9029461816957, -15.0141476304264, -16.74224131871, 
    -18.2676717222706, -19.7032882903104, -21.1346569643132, 
    -22.6435261325828, -24.3274544579203, -26.3282199110804, 
    -28.8866571762997, -32.4728171499292, -38.0393904829566, -27.6953287358666 ;

 aacgm_gm_lats =
  86.1408110343443, 75.8208444428181, 68.8217316552352, 60.063124351646, 
    50.6508693255777, 41.2874536006825, 32.2372769775103, 23.5912532699401, 
    15.5397401676606, 8.5731100054337, -7.10660016330614, -13.8991323763459, 
    -22.6091072092224, -31.720288799822, -41.2878618816532, 
    -51.5496830206068, -63.0200186762859, -70.1210442729992,
  83.9774633702212, 79.4584504860709, 73.1232062465901, 64.7366519590596, 
    55.6453807329812, 46.2743677172354, 36.7056549949636, 26.8242966368924, 
    16.845239972135, 8.18517497670915, -8.16589299185514, -16.2877724335302, 
    -25.4965317445022, -34.9270888212698, -44.7206644534399, 
    -55.1843821885905, -66.8518117245303, -69.5146024967299 ;

 aacgm_gm_lons =
  -151.839645671685, 80.032873562334, 51.5686003910971, 38.2527965556137, 
    30.6298617961532, 25.3061933272414, 20.7037991903455, 16.0662847165978, 
    11.3301650481058, 6.94085296657532, 3.3830960879891, 0.821603628248361, 
    -0.919868566303697, -2.21173093903996, -3.53251775368713, 
    -5.50368870993288, -8.94619308468165, 25.6785641609297,
  -145.218142931523, 57.6383740589023, 21.5417823925025, 6.49707224492552, 
    -1.91426752948519, -7.71611189526895, -12.1384952543716, 
    -15.4877766703428, -17.8004299420977, -19.231202542292, 
    -20.0585423333945, -20.4822840204513, -20.6161275402388, 
    -20.6478686116816, -20.8246751578698, -21.2593937438184, 
    -21.2343163068604, 19.9088658190448 ;
}
